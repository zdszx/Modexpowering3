module GroupPGLogic ( P_0_0,G_0_0,P_1_1,G_1_1,P_2_2,G_2_2,P_3_3,G_3_3,P_4_4,G_4_4,P_5_5,G_5_5,P_6_6,G_6_6,P_7_7,G_7_7,P_8_8,G_8_8,P_9_9,G_9_9,P_10_10,G_10_10,P_11_11,G_11_11,P_12_12,G_12_12,P_13_13,G_13_13,P_14_14,G_14_14,P_15_15,G_15_15,P_16_16,G_16_16,P_17_17,G_17_17,P_18_18,G_18_18,P_19_19,G_19_19,P_20_20,G_20_20,P_21_21,G_21_21,P_22_22,G_22_22,P_23_23,G_23_23,P_24_24,G_24_24,P_25_25,G_25_25,P_26_26,G_26_26,P_27_27,G_27_27,P_28_28,G_28_28,P_29_29,G_29_29,P_30_30,G_30_30,P_31_31,G_31_31,P_32_32,G_32_32,P_33_33,G_33_33,P_34_34,G_34_34,P_35_35,G_35_35,P_36_36,G_36_36,P_37_37,G_37_37,P_38_38,G_38_38,P_39_39,G_39_39,P_40_40,G_40_40,P_41_41,G_41_41,P_42_42,G_42_42,P_43_43,G_43_43,P_44_44,G_44_44,P_45_45,G_45_45,P_46_46,G_46_46,P_47_47,G_47_47,P_48_48,G_48_48,P_49_49,G_49_49,P_50_50,G_50_50,P_51_51,G_51_51,P_52_52,G_52_52,P_53_53,G_53_53,P_54_54,G_54_54,P_55_55,G_55_55,P_56_56,G_56_56,P_57_57,G_57_57,P_58_58,G_58_58,P_59_59,G_59_59,P_60_60,G_60_60,P_61_61,G_61_61,P_62_62,G_62_62,P_63_63,G_63_63,P_64_64,G_64_64,_P_0_0,_G_0_0,P_1_0,G_1_0,P_2_0,G_2_0,P_3_0,G_3_0,P_4_0,G_4_0,P_5_0,G_5_0,P_6_0,G_6_0,P_7_0,G_7_0,P_8_0,G_8_0,P_9_0,G_9_0,P_10_0,G_10_0,P_11_0,G_11_0,P_12_0,G_12_0,P_13_0,G_13_0,P_14_0,G_14_0,P_15_0,G_15_0,P_16_0,G_16_0,P_17_0,G_17_0,P_18_0,G_18_0,P_19_0,G_19_0,P_20_0,G_20_0,P_21_0,G_21_0,P_22_0,G_22_0,P_23_0,G_23_0,P_24_0,G_24_0,P_25_0,G_25_0,P_26_0,G_26_0,P_27_0,G_27_0,P_28_0,G_28_0,P_29_0,G_29_0,P_30_0,G_30_0,P_31_0,G_31_0,P_32_0,G_32_0,P_33_0,G_33_0,P_34_0,G_34_0,P_35_0,G_35_0,P_36_0,G_36_0,P_37_0,G_37_0,P_38_0,G_38_0,P_39_0,G_39_0,P_40_0,G_40_0,P_41_0,G_41_0,P_42_0,G_42_0,P_43_0,G_43_0,P_44_0,G_44_0,P_45_0,G_45_0,P_46_0,G_46_0,P_47_0,G_47_0,P_48_0,G_48_0,P_49_0,G_49_0,P_50_0,G_50_0,P_51_0,G_51_0,P_52_0,G_52_0,P_53_0,G_53_0,P_54_0,G_54_0,P_55_0,G_55_0,P_56_0,G_56_0,P_57_0,G_57_0,P_58_0,G_58_0,P_59_0,G_59_0,P_60_0,G_60_0,P_61_0,G_61_0,P_62_0,G_62_0,P_63_0,G_63_0,P_64_0,G_64_0 );
input P_0_0;
input G_0_0;
input P_1_1;
input G_1_1;
input P_2_2;
input G_2_2;
input P_3_3;
input G_3_3;
input P_4_4;
input G_4_4;
input P_5_5;
input G_5_5;
input P_6_6;
input G_6_6;
input P_7_7;
input G_7_7;
input P_8_8;
input G_8_8;
input P_9_9;
input G_9_9;
input P_10_10;
input G_10_10;
input P_11_11;
input G_11_11;
input P_12_12;
input G_12_12;
input P_13_13;
input G_13_13;
input P_14_14;
input G_14_14;
input P_15_15;
input G_15_15;
input P_16_16;
input G_16_16;
input P_17_17;
input G_17_17;
input P_18_18;
input G_18_18;
input P_19_19;
input G_19_19;
input P_20_20;
input G_20_20;
input P_21_21;
input G_21_21;
input P_22_22;
input G_22_22;
input P_23_23;
input G_23_23;
input P_24_24;
input G_24_24;
input P_25_25;
input G_25_25;
input P_26_26;
input G_26_26;
input P_27_27;
input G_27_27;
input P_28_28;
input G_28_28;
input P_29_29;
input G_29_29;
input P_30_30;
input G_30_30;
input P_31_31;
input G_31_31;
input P_32_32;
input G_32_32;
input P_33_33;
input G_33_33;
input P_34_34;
input G_34_34;
input P_35_35;
input G_35_35;
input P_36_36;
input G_36_36;
input P_37_37;
input G_37_37;
input P_38_38;
input G_38_38;
input P_39_39;
input G_39_39;
input P_40_40;
input G_40_40;
input P_41_41;
input G_41_41;
input P_42_42;
input G_42_42;
input P_43_43;
input G_43_43;
input P_44_44;
input G_44_44;
input P_45_45;
input G_45_45;
input P_46_46;
input G_46_46;
input P_47_47;
input G_47_47;
input P_48_48;
input G_48_48;
input P_49_49;
input G_49_49;
input P_50_50;
input G_50_50;
input P_51_51;
input G_51_51;
input P_52_52;
input G_52_52;
input P_53_53;
input G_53_53;
input P_54_54;
input G_54_54;
input P_55_55;
input G_55_55;
input P_56_56;
input G_56_56;
input P_57_57;
input G_57_57;
input P_58_58;
input G_58_58;
input P_59_59;
input G_59_59;
input P_60_60;
input G_60_60;
input P_61_61;
input G_61_61;
input P_62_62;
input G_62_62;
input P_63_63;
input G_63_63;
input P_64_64;
input G_64_64;
output _P_0_0;
output _G_0_0;
output P_1_0;
output G_1_0;
output P_2_0;
output G_2_0;
output P_3_0;
output G_3_0;
output P_4_0;
output G_4_0;
output P_5_0;
output G_5_0;
output P_6_0;
output G_6_0;
output P_7_0;
output G_7_0;
output P_8_0;
output G_8_0;
output P_9_0;
output G_9_0;
output P_10_0;
output G_10_0;
output P_11_0;
output G_11_0;
output P_12_0;
output G_12_0;
output P_13_0;
output G_13_0;
output P_14_0;
output G_14_0;
output P_15_0;
output G_15_0;
output P_16_0;
output G_16_0;
output P_17_0;
output G_17_0;
output P_18_0;
output G_18_0;
output P_19_0;
output G_19_0;
output P_20_0;
output G_20_0;
output P_21_0;
output G_21_0;
output P_22_0;
output G_22_0;
output P_23_0;
output G_23_0;
output P_24_0;
output G_24_0;
output P_25_0;
output G_25_0;
output P_26_0;
output G_26_0;
output P_27_0;
output G_27_0;
output P_28_0;
output G_28_0;
output P_29_0;
output G_29_0;
output P_30_0;
output G_30_0;
output P_31_0;
output G_31_0;
output P_32_0;
output G_32_0;
output P_33_0;
output G_33_0;
output P_34_0;
output G_34_0;
output P_35_0;
output G_35_0;
output P_36_0;
output G_36_0;
output P_37_0;
output G_37_0;
output P_38_0;
output G_38_0;
output P_39_0;
output G_39_0;
output P_40_0;
output G_40_0;
output P_41_0;
output G_41_0;
output P_42_0;
output G_42_0;
output P_43_0;
output G_43_0;
output P_44_0;
output G_44_0;
output P_45_0;
output G_45_0;
output P_46_0;
output G_46_0;
output P_47_0;
output G_47_0;
output P_48_0;
output G_48_0;
output P_49_0;
output G_49_0;
output P_50_0;
output G_50_0;
output P_51_0;
output G_51_0;
output P_52_0;
output G_52_0;
output P_53_0;
output G_53_0;
output P_54_0;
output G_54_0;
output P_55_0;
output G_55_0;
output P_56_0;
output G_56_0;
output P_57_0;
output G_57_0;
output P_58_0;
output G_58_0;
output P_59_0;
output G_59_0;
output P_60_0;
output G_60_0;
output P_61_0;
output G_61_0;
output P_62_0;
output G_62_0;
output P_63_0;
output G_63_0;
output P_64_0;
output G_64_0;
wire G_3_2;
wire P_3_2;
wire G_5_4;
wire P_5_4;
wire G_7_6;
wire P_7_6;
wire G_9_8;
wire P_9_8;
wire G_11_10;
wire P_11_10;
wire G_13_12;
wire P_13_12;
wire G_15_14;
wire P_15_14;
wire G_17_16;
wire P_17_16;
wire G_19_18;
wire P_19_18;
wire G_21_20;
wire P_21_20;
wire G_23_22;
wire P_23_22;
wire G_25_24;
wire P_25_24;
wire G_27_26;
wire P_27_26;
wire G_29_28;
wire P_29_28;
wire G_31_30;
wire P_31_30;
wire G_33_32;
wire P_33_32;
wire G_35_34;
wire P_35_34;
wire G_37_36;
wire P_37_36;
wire G_39_38;
wire P_39_38;
wire G_41_40;
wire P_41_40;
wire G_43_42;
wire P_43_42;
wire G_45_44;
wire P_45_44;
wire G_47_46;
wire P_47_46;
wire G_49_48;
wire P_49_48;
wire G_51_50;
wire P_51_50;
wire G_53_52;
wire P_53_52;
wire G_55_54;
wire P_55_54;
wire G_57_56;
wire P_57_56;
wire G_59_58;
wire P_59_58;
wire G_61_60;
wire P_61_60;
wire G_63_62;
wire P_63_62;
wire G_7_4;
wire P_7_4;
wire G_11_8;
wire P_11_8;
wire G_15_12;
wire P_15_12;
wire G_19_16;
wire P_19_16;
wire G_23_20;
wire P_23_20;
wire G_27_24;
wire P_27_24;
wire G_31_28;
wire P_31_28;
wire G_35_32;
wire P_35_32;
wire G_39_36;
wire P_39_36;
wire G_43_40;
wire P_43_40;
wire G_47_44;
wire P_47_44;
wire G_51_48;
wire P_51_48;
wire G_55_52;
wire P_55_52;
wire G_59_56;
wire P_59_56;
wire G_63_60;
wire P_63_60;
wire G_15_8;
wire P_15_8;
wire G_23_16;
wire P_23_16;
wire G_31_24;
wire P_31_24;
wire G_39_32;
wire P_39_32;
wire G_47_40;
wire P_47_40;
wire G_55_48;
wire P_55_48;
wire G_63_56;
wire P_63_56;
wire G_31_16;
wire P_31_16;
wire G_47_32;
wire P_47_32;
wire G_63_48;
wire P_63_48;
wire G_63_32;
wire P_63_32;
GrayBlock gray_block_1_0(.G_i_k(G_1_1),.P_i_k(P_1_1),.G_km1_j(G_0_0),.G_i_j(G_1_0));
BlackBlock black_block_3_2(.G_i_k(G_3_3),.P_i_k(P_3_3),.G_km1_j(G_2_2),.P_km1_j(P_2_2),.G_i_j(G_3_2),.P_i_j(P_3_2));
BlackBlock black_block_5_4(.G_i_k(G_5_5),.P_i_k(P_5_5),.G_km1_j(G_4_4),.P_km1_j(P_4_4),.G_i_j(G_5_4),.P_i_j(P_5_4));
BlackBlock black_block_7_6(.G_i_k(G_7_7),.P_i_k(P_7_7),.G_km1_j(G_6_6),.P_km1_j(P_6_6),.G_i_j(G_7_6),.P_i_j(P_7_6));
BlackBlock black_block_9_8(.G_i_k(G_9_9),.P_i_k(P_9_9),.G_km1_j(G_8_8),.P_km1_j(P_8_8),.G_i_j(G_9_8),.P_i_j(P_9_8));
BlackBlock black_block_11_10(.G_i_k(G_11_11),.P_i_k(P_11_11),.G_km1_j(G_10_10),.P_km1_j(P_10_10),.G_i_j(G_11_10),.P_i_j(P_11_10));
BlackBlock black_block_13_12(.G_i_k(G_13_13),.P_i_k(P_13_13),.G_km1_j(G_12_12),.P_km1_j(P_12_12),.G_i_j(G_13_12),.P_i_j(P_13_12));
BlackBlock black_block_15_14(.G_i_k(G_15_15),.P_i_k(P_15_15),.G_km1_j(G_14_14),.P_km1_j(P_14_14),.G_i_j(G_15_14),.P_i_j(P_15_14));
BlackBlock black_block_17_16(.G_i_k(G_17_17),.P_i_k(P_17_17),.G_km1_j(G_16_16),.P_km1_j(P_16_16),.G_i_j(G_17_16),.P_i_j(P_17_16));
BlackBlock black_block_19_18(.G_i_k(G_19_19),.P_i_k(P_19_19),.G_km1_j(G_18_18),.P_km1_j(P_18_18),.G_i_j(G_19_18),.P_i_j(P_19_18));
BlackBlock black_block_21_20(.G_i_k(G_21_21),.P_i_k(P_21_21),.G_km1_j(G_20_20),.P_km1_j(P_20_20),.G_i_j(G_21_20),.P_i_j(P_21_20));
BlackBlock black_block_23_22(.G_i_k(G_23_23),.P_i_k(P_23_23),.G_km1_j(G_22_22),.P_km1_j(P_22_22),.G_i_j(G_23_22),.P_i_j(P_23_22));
BlackBlock black_block_25_24(.G_i_k(G_25_25),.P_i_k(P_25_25),.G_km1_j(G_24_24),.P_km1_j(P_24_24),.G_i_j(G_25_24),.P_i_j(P_25_24));
BlackBlock black_block_27_26(.G_i_k(G_27_27),.P_i_k(P_27_27),.G_km1_j(G_26_26),.P_km1_j(P_26_26),.G_i_j(G_27_26),.P_i_j(P_27_26));
BlackBlock black_block_29_28(.G_i_k(G_29_29),.P_i_k(P_29_29),.G_km1_j(G_28_28),.P_km1_j(P_28_28),.G_i_j(G_29_28),.P_i_j(P_29_28));
BlackBlock black_block_31_30(.G_i_k(G_31_31),.P_i_k(P_31_31),.G_km1_j(G_30_30),.P_km1_j(P_30_30),.G_i_j(G_31_30),.P_i_j(P_31_30));
BlackBlock black_block_33_32(.G_i_k(G_33_33),.P_i_k(P_33_33),.G_km1_j(G_32_32),.P_km1_j(P_32_32),.G_i_j(G_33_32),.P_i_j(P_33_32));
BlackBlock black_block_35_34(.G_i_k(G_35_35),.P_i_k(P_35_35),.G_km1_j(G_34_34),.P_km1_j(P_34_34),.G_i_j(G_35_34),.P_i_j(P_35_34));
BlackBlock black_block_37_36(.G_i_k(G_37_37),.P_i_k(P_37_37),.G_km1_j(G_36_36),.P_km1_j(P_36_36),.G_i_j(G_37_36),.P_i_j(P_37_36));
BlackBlock black_block_39_38(.G_i_k(G_39_39),.P_i_k(P_39_39),.G_km1_j(G_38_38),.P_km1_j(P_38_38),.G_i_j(G_39_38),.P_i_j(P_39_38));
BlackBlock black_block_41_40(.G_i_k(G_41_41),.P_i_k(P_41_41),.G_km1_j(G_40_40),.P_km1_j(P_40_40),.G_i_j(G_41_40),.P_i_j(P_41_40));
BlackBlock black_block_43_42(.G_i_k(G_43_43),.P_i_k(P_43_43),.G_km1_j(G_42_42),.P_km1_j(P_42_42),.G_i_j(G_43_42),.P_i_j(P_43_42));
BlackBlock black_block_45_44(.G_i_k(G_45_45),.P_i_k(P_45_45),.G_km1_j(G_44_44),.P_km1_j(P_44_44),.G_i_j(G_45_44),.P_i_j(P_45_44));
BlackBlock black_block_47_46(.G_i_k(G_47_47),.P_i_k(P_47_47),.G_km1_j(G_46_46),.P_km1_j(P_46_46),.G_i_j(G_47_46),.P_i_j(P_47_46));
BlackBlock black_block_49_48(.G_i_k(G_49_49),.P_i_k(P_49_49),.G_km1_j(G_48_48),.P_km1_j(P_48_48),.G_i_j(G_49_48),.P_i_j(P_49_48));
BlackBlock black_block_51_50(.G_i_k(G_51_51),.P_i_k(P_51_51),.G_km1_j(G_50_50),.P_km1_j(P_50_50),.G_i_j(G_51_50),.P_i_j(P_51_50));
BlackBlock black_block_53_52(.G_i_k(G_53_53),.P_i_k(P_53_53),.G_km1_j(G_52_52),.P_km1_j(P_52_52),.G_i_j(G_53_52),.P_i_j(P_53_52));
BlackBlock black_block_55_54(.G_i_k(G_55_55),.P_i_k(P_55_55),.G_km1_j(G_54_54),.P_km1_j(P_54_54),.G_i_j(G_55_54),.P_i_j(P_55_54));
BlackBlock black_block_57_56(.G_i_k(G_57_57),.P_i_k(P_57_57),.G_km1_j(G_56_56),.P_km1_j(P_56_56),.G_i_j(G_57_56),.P_i_j(P_57_56));
BlackBlock black_block_59_58(.G_i_k(G_59_59),.P_i_k(P_59_59),.G_km1_j(G_58_58),.P_km1_j(P_58_58),.G_i_j(G_59_58),.P_i_j(P_59_58));
BlackBlock black_block_61_60(.G_i_k(G_61_61),.P_i_k(P_61_61),.G_km1_j(G_60_60),.P_km1_j(P_60_60),.G_i_j(G_61_60),.P_i_j(P_61_60));
BlackBlock black_block_63_62(.G_i_k(G_63_63),.P_i_k(P_63_63),.G_km1_j(G_62_62),.P_km1_j(P_62_62),.G_i_j(G_63_62),.P_i_j(P_63_62));
GrayBlock gray_block_3_0(.G_i_k(G_3_2),.P_i_k(P_3_2),.G_km1_j(G_1_0),.G_i_j(G_3_0));
BlackBlock black_block_7_4(.G_i_k(G_7_6),.P_i_k(P_7_6),.G_km1_j(G_5_4),.P_km1_j(P_5_4),.G_i_j(G_7_4),.P_i_j(P_7_4));
BlackBlock black_block_11_8(.G_i_k(G_11_10),.P_i_k(P_11_10),.G_km1_j(G_9_8),.P_km1_j(P_9_8),.G_i_j(G_11_8),.P_i_j(P_11_8));
BlackBlock black_block_15_12(.G_i_k(G_15_14),.P_i_k(P_15_14),.G_km1_j(G_13_12),.P_km1_j(P_13_12),.G_i_j(G_15_12),.P_i_j(P_15_12));
BlackBlock black_block_19_16(.G_i_k(G_19_18),.P_i_k(P_19_18),.G_km1_j(G_17_16),.P_km1_j(P_17_16),.G_i_j(G_19_16),.P_i_j(P_19_16));
BlackBlock black_block_23_20(.G_i_k(G_23_22),.P_i_k(P_23_22),.G_km1_j(G_21_20),.P_km1_j(P_21_20),.G_i_j(G_23_20),.P_i_j(P_23_20));
BlackBlock black_block_27_24(.G_i_k(G_27_26),.P_i_k(P_27_26),.G_km1_j(G_25_24),.P_km1_j(P_25_24),.G_i_j(G_27_24),.P_i_j(P_27_24));
BlackBlock black_block_31_28(.G_i_k(G_31_30),.P_i_k(P_31_30),.G_km1_j(G_29_28),.P_km1_j(P_29_28),.G_i_j(G_31_28),.P_i_j(P_31_28));
BlackBlock black_block_35_32(.G_i_k(G_35_34),.P_i_k(P_35_34),.G_km1_j(G_33_32),.P_km1_j(P_33_32),.G_i_j(G_35_32),.P_i_j(P_35_32));
BlackBlock black_block_39_36(.G_i_k(G_39_38),.P_i_k(P_39_38),.G_km1_j(G_37_36),.P_km1_j(P_37_36),.G_i_j(G_39_36),.P_i_j(P_39_36));
BlackBlock black_block_43_40(.G_i_k(G_43_42),.P_i_k(P_43_42),.G_km1_j(G_41_40),.P_km1_j(P_41_40),.G_i_j(G_43_40),.P_i_j(P_43_40));
BlackBlock black_block_47_44(.G_i_k(G_47_46),.P_i_k(P_47_46),.G_km1_j(G_45_44),.P_km1_j(P_45_44),.G_i_j(G_47_44),.P_i_j(P_47_44));
BlackBlock black_block_51_48(.G_i_k(G_51_50),.P_i_k(P_51_50),.G_km1_j(G_49_48),.P_km1_j(P_49_48),.G_i_j(G_51_48),.P_i_j(P_51_48));
BlackBlock black_block_55_52(.G_i_k(G_55_54),.P_i_k(P_55_54),.G_km1_j(G_53_52),.P_km1_j(P_53_52),.G_i_j(G_55_52),.P_i_j(P_55_52));
BlackBlock black_block_59_56(.G_i_k(G_59_58),.P_i_k(P_59_58),.G_km1_j(G_57_56),.P_km1_j(P_57_56),.G_i_j(G_59_56),.P_i_j(P_59_56));
BlackBlock black_block_63_60(.G_i_k(G_63_62),.P_i_k(P_63_62),.G_km1_j(G_61_60),.P_km1_j(P_61_60),.G_i_j(G_63_60),.P_i_j(P_63_60));
GrayBlock gray_block_7_0(.G_i_k(G_7_4),.P_i_k(P_7_4),.G_km1_j(G_3_0),.G_i_j(G_7_0));
BlackBlock black_block_15_8(.G_i_k(G_15_12),.P_i_k(P_15_12),.G_km1_j(G_11_8),.P_km1_j(P_11_8),.G_i_j(G_15_8),.P_i_j(P_15_8));
BlackBlock black_block_23_16(.G_i_k(G_23_20),.P_i_k(P_23_20),.G_km1_j(G_19_16),.P_km1_j(P_19_16),.G_i_j(G_23_16),.P_i_j(P_23_16));
BlackBlock black_block_31_24(.G_i_k(G_31_28),.P_i_k(P_31_28),.G_km1_j(G_27_24),.P_km1_j(P_27_24),.G_i_j(G_31_24),.P_i_j(P_31_24));
BlackBlock black_block_39_32(.G_i_k(G_39_36),.P_i_k(P_39_36),.G_km1_j(G_35_32),.P_km1_j(P_35_32),.G_i_j(G_39_32),.P_i_j(P_39_32));
BlackBlock black_block_47_40(.G_i_k(G_47_44),.P_i_k(P_47_44),.G_km1_j(G_43_40),.P_km1_j(P_43_40),.G_i_j(G_47_40),.P_i_j(P_47_40));
BlackBlock black_block_55_48(.G_i_k(G_55_52),.P_i_k(P_55_52),.G_km1_j(G_51_48),.P_km1_j(P_51_48),.G_i_j(G_55_48),.P_i_j(P_55_48));
BlackBlock black_block_63_56(.G_i_k(G_63_60),.P_i_k(P_63_60),.G_km1_j(G_59_56),.P_km1_j(P_59_56),.G_i_j(G_63_56),.P_i_j(P_63_56));
GrayBlock gray_block_15_0(.G_i_k(G_15_8),.P_i_k(P_15_8),.G_km1_j(G_7_0),.G_i_j(G_15_0));
BlackBlock black_block_31_16(.G_i_k(G_31_24),.P_i_k(P_31_24),.G_km1_j(G_23_16),.P_km1_j(P_23_16),.G_i_j(G_31_16),.P_i_j(P_31_16));
BlackBlock black_block_47_32(.G_i_k(G_47_40),.P_i_k(P_47_40),.G_km1_j(G_39_32),.P_km1_j(P_39_32),.G_i_j(G_47_32),.P_i_j(P_47_32));
BlackBlock black_block_63_48(.G_i_k(G_63_56),.P_i_k(P_63_56),.G_km1_j(G_55_48),.P_km1_j(P_55_48),.G_i_j(G_63_48),.P_i_j(P_63_48));
GrayBlock gray_block_31_0(.G_i_k(G_31_16),.P_i_k(P_31_16),.G_km1_j(G_15_0),.G_i_j(G_31_0));
BlackBlock black_block_63_32(.G_i_k(G_63_48),.P_i_k(P_63_48),.G_km1_j(G_47_32),.P_km1_j(P_47_32),.G_i_j(G_63_32),.P_i_j(P_63_32));
GrayBlock gray_block_63_0(.G_i_k(G_63_32),.P_i_k(P_63_32),.G_km1_j(G_31_0),.G_i_j(G_63_0));
GrayBlock gray_block_47_31(.G_i_k(G_47_32),.P_i_k(P_47_32),.G_km1_j(G_31_0),.G_i_j(G_47_0));
GrayBlock gray_block_23_15(.G_i_k(G_23_16),.P_i_k(P_23_16),.G_km1_j(G_15_0),.G_i_j(G_23_0));
GrayBlock gray_block_39_31(.G_i_k(G_39_32),.P_i_k(P_39_32),.G_km1_j(G_31_0),.G_i_j(G_39_0));
GrayBlock gray_block_55_47(.G_i_k(G_55_48),.P_i_k(P_55_48),.G_km1_j(G_47_0),.G_i_j(G_55_0));
GrayBlock gray_block_11_7(.G_i_k(G_11_8),.P_i_k(P_11_8),.G_km1_j(G_7_0),.G_i_j(G_11_0));
GrayBlock gray_block_19_15(.G_i_k(G_19_16),.P_i_k(P_19_16),.G_km1_j(G_15_0),.G_i_j(G_19_0));
GrayBlock gray_block_27_23(.G_i_k(G_27_24),.P_i_k(P_27_24),.G_km1_j(G_23_0),.G_i_j(G_27_0));
GrayBlock gray_block_35_31(.G_i_k(G_35_32),.P_i_k(P_35_32),.G_km1_j(G_31_0),.G_i_j(G_35_0));
GrayBlock gray_block_43_39(.G_i_k(G_43_40),.P_i_k(P_43_40),.G_km1_j(G_39_0),.G_i_j(G_43_0));
GrayBlock gray_block_51_47(.G_i_k(G_51_48),.P_i_k(P_51_48),.G_km1_j(G_47_0),.G_i_j(G_51_0));
GrayBlock gray_block_59_55(.G_i_k(G_59_56),.P_i_k(P_59_56),.G_km1_j(G_55_0),.G_i_j(G_59_0));
GrayBlock gray_block_5_3(.G_i_k(G_5_4),.P_i_k(P_5_4),.G_km1_j(G_3_0),.G_i_j(G_5_0));
GrayBlock gray_block_9_7(.G_i_k(G_9_8),.P_i_k(P_9_8),.G_km1_j(G_7_0),.G_i_j(G_9_0));
GrayBlock gray_block_13_11(.G_i_k(G_13_12),.P_i_k(P_13_12),.G_km1_j(G_11_0),.G_i_j(G_13_0));
GrayBlock gray_block_17_15(.G_i_k(G_17_16),.P_i_k(P_17_16),.G_km1_j(G_15_0),.G_i_j(G_17_0));
GrayBlock gray_block_21_19(.G_i_k(G_21_20),.P_i_k(P_21_20),.G_km1_j(G_19_0),.G_i_j(G_21_0));
GrayBlock gray_block_25_23(.G_i_k(G_25_24),.P_i_k(P_25_24),.G_km1_j(G_23_0),.G_i_j(G_25_0));
GrayBlock gray_block_29_27(.G_i_k(G_29_28),.P_i_k(P_29_28),.G_km1_j(G_27_0),.G_i_j(G_29_0));
GrayBlock gray_block_33_31(.G_i_k(G_33_32),.P_i_k(P_33_32),.G_km1_j(G_31_0),.G_i_j(G_33_0));
GrayBlock gray_block_37_35(.G_i_k(G_37_36),.P_i_k(P_37_36),.G_km1_j(G_35_0),.G_i_j(G_37_0));
GrayBlock gray_block_41_39(.G_i_k(G_41_40),.P_i_k(P_41_40),.G_km1_j(G_39_0),.G_i_j(G_41_0));
GrayBlock gray_block_45_43(.G_i_k(G_45_44),.P_i_k(P_45_44),.G_km1_j(G_43_0),.G_i_j(G_45_0));
GrayBlock gray_block_49_47(.G_i_k(G_49_48),.P_i_k(P_49_48),.G_km1_j(G_47_0),.G_i_j(G_49_0));
GrayBlock gray_block_53_51(.G_i_k(G_53_52),.P_i_k(P_53_52),.G_km1_j(G_51_0),.G_i_j(G_53_0));
GrayBlock gray_block_57_55(.G_i_k(G_57_56),.P_i_k(P_57_56),.G_km1_j(G_55_0),.G_i_j(G_57_0));
GrayBlock gray_block_61_59(.G_i_k(G_61_60),.P_i_k(P_61_60),.G_km1_j(G_59_0),.G_i_j(G_61_0));
GrayBlock gray_block_2_1(.G_i_k(G_2_2),.P_i_k(P_2_2),.G_km1_j(G_1_0),.G_i_j(G_2_0));
GrayBlock gray_block_4_3(.G_i_k(G_4_4),.P_i_k(P_4_4),.G_km1_j(G_3_0),.G_i_j(G_4_0));
GrayBlock gray_block_6_5(.G_i_k(G_6_6),.P_i_k(P_6_6),.G_km1_j(G_5_0),.G_i_j(G_6_0));
GrayBlock gray_block_8_7(.G_i_k(G_8_8),.P_i_k(P_8_8),.G_km1_j(G_7_0),.G_i_j(G_8_0));
GrayBlock gray_block_10_9(.G_i_k(G_10_10),.P_i_k(P_10_10),.G_km1_j(G_9_0),.G_i_j(G_10_0));
GrayBlock gray_block_12_11(.G_i_k(G_12_12),.P_i_k(P_12_12),.G_km1_j(G_11_0),.G_i_j(G_12_0));
GrayBlock gray_block_14_13(.G_i_k(G_14_14),.P_i_k(P_14_14),.G_km1_j(G_13_0),.G_i_j(G_14_0));
GrayBlock gray_block_16_15(.G_i_k(G_16_16),.P_i_k(P_16_16),.G_km1_j(G_15_0),.G_i_j(G_16_0));
GrayBlock gray_block_18_17(.G_i_k(G_18_18),.P_i_k(P_18_18),.G_km1_j(G_17_0),.G_i_j(G_18_0));
GrayBlock gray_block_20_19(.G_i_k(G_20_20),.P_i_k(P_20_20),.G_km1_j(G_19_0),.G_i_j(G_20_0));
GrayBlock gray_block_22_21(.G_i_k(G_22_22),.P_i_k(P_22_22),.G_km1_j(G_21_0),.G_i_j(G_22_0));
GrayBlock gray_block_24_23(.G_i_k(G_24_24),.P_i_k(P_24_24),.G_km1_j(G_23_0),.G_i_j(G_24_0));
GrayBlock gray_block_26_25(.G_i_k(G_26_26),.P_i_k(P_26_26),.G_km1_j(G_25_0),.G_i_j(G_26_0));
GrayBlock gray_block_28_27(.G_i_k(G_28_28),.P_i_k(P_28_28),.G_km1_j(G_27_0),.G_i_j(G_28_0));
GrayBlock gray_block_30_29(.G_i_k(G_30_30),.P_i_k(P_30_30),.G_km1_j(G_29_0),.G_i_j(G_30_0));
GrayBlock gray_block_32_31(.G_i_k(G_32_32),.P_i_k(P_32_32),.G_km1_j(G_31_0),.G_i_j(G_32_0));
GrayBlock gray_block_34_33(.G_i_k(G_34_34),.P_i_k(P_34_34),.G_km1_j(G_33_0),.G_i_j(G_34_0));
GrayBlock gray_block_36_35(.G_i_k(G_36_36),.P_i_k(P_36_36),.G_km1_j(G_35_0),.G_i_j(G_36_0));
GrayBlock gray_block_38_37(.G_i_k(G_38_38),.P_i_k(P_38_38),.G_km1_j(G_37_0),.G_i_j(G_38_0));
GrayBlock gray_block_40_39(.G_i_k(G_40_40),.P_i_k(P_40_40),.G_km1_j(G_39_0),.G_i_j(G_40_0));
GrayBlock gray_block_42_41(.G_i_k(G_42_42),.P_i_k(P_42_42),.G_km1_j(G_41_0),.G_i_j(G_42_0));
GrayBlock gray_block_44_43(.G_i_k(G_44_44),.P_i_k(P_44_44),.G_km1_j(G_43_0),.G_i_j(G_44_0));
GrayBlock gray_block_46_45(.G_i_k(G_46_46),.P_i_k(P_46_46),.G_km1_j(G_45_0),.G_i_j(G_46_0));
GrayBlock gray_block_48_47(.G_i_k(G_48_48),.P_i_k(P_48_48),.G_km1_j(G_47_0),.G_i_j(G_48_0));
GrayBlock gray_block_50_49(.G_i_k(G_50_50),.P_i_k(P_50_50),.G_km1_j(G_49_0),.G_i_j(G_50_0));
GrayBlock gray_block_52_51(.G_i_k(G_52_52),.P_i_k(P_52_52),.G_km1_j(G_51_0),.G_i_j(G_52_0));
GrayBlock gray_block_54_53(.G_i_k(G_54_54),.P_i_k(P_54_54),.G_km1_j(G_53_0),.G_i_j(G_54_0));
GrayBlock gray_block_56_55(.G_i_k(G_56_56),.P_i_k(P_56_56),.G_km1_j(G_55_0),.G_i_j(G_56_0));
GrayBlock gray_block_58_57(.G_i_k(G_58_58),.P_i_k(P_58_58),.G_km1_j(G_57_0),.G_i_j(G_58_0));
GrayBlock gray_block_60_59(.G_i_k(G_60_60),.P_i_k(P_60_60),.G_km1_j(G_59_0),.G_i_j(G_60_0));
GrayBlock gray_block_62_61(.G_i_k(G_62_62),.P_i_k(P_62_62),.G_km1_j(G_61_0),.G_i_j(G_62_0));
GrayBlock gray_block_64_63(.G_i_k(G_64_64),.P_i_k(P_64_64),.G_km1_j(G_63_0),.G_i_j(G_64_0));
assign _P_0_0 = P_0_0 ;
assign _G_0_0 = G_0_0 ;
endmodule
