module GroupPGLogic ( P_0_0,G_0_0,P_1_1,G_1_1,P_2_2,G_2_2,P_3_3,G_3_3,P_4_4,G_4_4,P_5_5,G_5_5,P_6_6,G_6_6,P_7_7,G_7_7,P_8_8,G_8_8,P_9_9,G_9_9,P_10_10,G_10_10,P_11_11,G_11_11,P_12_12,G_12_12,P_13_13,G_13_13,P_14_14,G_14_14,P_15_15,G_15_15,P_16_16,G_16_16,P_17_17,G_17_17,P_18_18,G_18_18,P_19_19,G_19_19,P_20_20,G_20_20,P_21_21,G_21_21,P_22_22,G_22_22,P_23_23,G_23_23,P_24_24,G_24_24,P_25_25,G_25_25,P_26_26,G_26_26,P_27_27,G_27_27,P_28_28,G_28_28,P_29_29,G_29_29,P_30_30,G_30_30,P_31_31,G_31_31,P_32_32,G_32_32,_P_0_0,_G_0_0,P_1_0,G_1_0,P_2_0,G_2_0,P_3_0,G_3_0,P_4_0,G_4_0,P_5_0,G_5_0,P_6_0,G_6_0,P_7_0,G_7_0,P_8_0,G_8_0,P_9_0,G_9_0,P_10_0,G_10_0,P_11_0,G_11_0,P_12_0,G_12_0,P_13_0,G_13_0,P_14_0,G_14_0,P_15_0,G_15_0,P_16_0,G_16_0,P_17_0,G_17_0,P_18_0,G_18_0,P_19_0,G_19_0,P_20_0,G_20_0,P_21_0,G_21_0,P_22_0,G_22_0,P_23_0,G_23_0,P_24_0,G_24_0,P_25_0,G_25_0,P_26_0,G_26_0,P_27_0,G_27_0,P_28_0,G_28_0,P_29_0,G_29_0,P_30_0,G_30_0,P_31_0,G_31_0,P_32_0,G_32_0 );
input P_0_0;
input G_0_0;
input P_1_1;
input G_1_1;
input P_2_2;
input G_2_2;
input P_3_3;
input G_3_3;
input P_4_4;
input G_4_4;
input P_5_5;
input G_5_5;
input P_6_6;
input G_6_6;
input P_7_7;
input G_7_7;
input P_8_8;
input G_8_8;
input P_9_9;
input G_9_9;
input P_10_10;
input G_10_10;
input P_11_11;
input G_11_11;
input P_12_12;
input G_12_12;
input P_13_13;
input G_13_13;
input P_14_14;
input G_14_14;
input P_15_15;
input G_15_15;
input P_16_16;
input G_16_16;
input P_17_17;
input G_17_17;
input P_18_18;
input G_18_18;
input P_19_19;
input G_19_19;
input P_20_20;
input G_20_20;
input P_21_21;
input G_21_21;
input P_22_22;
input G_22_22;
input P_23_23;
input G_23_23;
input P_24_24;
input G_24_24;
input P_25_25;
input G_25_25;
input P_26_26;
input G_26_26;
input P_27_27;
input G_27_27;
input P_28_28;
input G_28_28;
input P_29_29;
input G_29_29;
input P_30_30;
input G_30_30;
input P_31_31;
input G_31_31;
input P_32_32;
input G_32_32;
output _P_0_0;
output _G_0_0;
output P_1_0;
output G_1_0;
output P_2_0;
output G_2_0;
output P_3_0;
output G_3_0;
output P_4_0;
output G_4_0;
output P_5_0;
output G_5_0;
output P_6_0;
output G_6_0;
output P_7_0;
output G_7_0;
output P_8_0;
output G_8_0;
output P_9_0;
output G_9_0;
output P_10_0;
output G_10_0;
output P_11_0;
output G_11_0;
output P_12_0;
output G_12_0;
output P_13_0;
output G_13_0;
output P_14_0;
output G_14_0;
output P_15_0;
output G_15_0;
output P_16_0;
output G_16_0;
output P_17_0;
output G_17_0;
output P_18_0;
output G_18_0;
output P_19_0;
output G_19_0;
output P_20_0;
output G_20_0;
output P_21_0;
output G_21_0;
output P_22_0;
output G_22_0;
output P_23_0;
output G_23_0;
output P_24_0;
output G_24_0;
output P_25_0;
output G_25_0;
output P_26_0;
output G_26_0;
output P_27_0;
output G_27_0;
output P_28_0;
output G_28_0;
output P_29_0;
output G_29_0;
output P_30_0;
output G_30_0;
output P_31_0;
output G_31_0;
output P_32_0;
output G_32_0;
wire G_3_2;
wire P_3_2;
wire G_5_4;
wire P_5_4;
wire G_7_6;
wire P_7_6;
wire G_9_8;
wire P_9_8;
wire G_11_10;
wire P_11_10;
wire G_13_12;
wire P_13_12;
wire G_15_14;
wire P_15_14;
wire G_17_16;
wire P_17_16;
wire G_19_18;
wire P_19_18;
wire G_21_20;
wire P_21_20;
wire G_23_22;
wire P_23_22;
wire G_25_24;
wire P_25_24;
wire G_27_26;
wire P_27_26;
wire G_29_28;
wire P_29_28;
wire G_31_30;
wire P_31_30;
wire G_7_4;
wire P_7_4;
wire G_11_8;
wire P_11_8;
wire G_15_12;
wire P_15_12;
wire G_19_16;
wire P_19_16;
wire G_23_20;
wire P_23_20;
wire G_27_24;
wire P_27_24;
wire G_31_28;
wire P_31_28;
wire G_15_8;
wire P_15_8;
wire G_23_16;
wire P_23_16;
wire G_31_24;
wire P_31_24;
wire G_31_16;
wire P_31_16;
GrayBlock gray_block_1_0(.G_i_k(G_1_1),.P_i_k(P_1_1),.G_km1_j(G_0_0),.G_i_j(G_1_0));
BlackBlock black_block_3_2(.G_i_k(G_3_3),.P_i_k(P_3_3),.G_km1_j(G_2_2),.P_km1_j(P_2_2),.G_i_j(G_3_2),.P_i_j(P_3_2));
BlackBlock black_block_5_4(.G_i_k(G_5_5),.P_i_k(P_5_5),.G_km1_j(G_4_4),.P_km1_j(P_4_4),.G_i_j(G_5_4),.P_i_j(P_5_4));
BlackBlock black_block_7_6(.G_i_k(G_7_7),.P_i_k(P_7_7),.G_km1_j(G_6_6),.P_km1_j(P_6_6),.G_i_j(G_7_6),.P_i_j(P_7_6));
BlackBlock black_block_9_8(.G_i_k(G_9_9),.P_i_k(P_9_9),.G_km1_j(G_8_8),.P_km1_j(P_8_8),.G_i_j(G_9_8),.P_i_j(P_9_8));
BlackBlock black_block_11_10(.G_i_k(G_11_11),.P_i_k(P_11_11),.G_km1_j(G_10_10),.P_km1_j(P_10_10),.G_i_j(G_11_10),.P_i_j(P_11_10));
BlackBlock black_block_13_12(.G_i_k(G_13_13),.P_i_k(P_13_13),.G_km1_j(G_12_12),.P_km1_j(P_12_12),.G_i_j(G_13_12),.P_i_j(P_13_12));
BlackBlock black_block_15_14(.G_i_k(G_15_15),.P_i_k(P_15_15),.G_km1_j(G_14_14),.P_km1_j(P_14_14),.G_i_j(G_15_14),.P_i_j(P_15_14));
BlackBlock black_block_17_16(.G_i_k(G_17_17),.P_i_k(P_17_17),.G_km1_j(G_16_16),.P_km1_j(P_16_16),.G_i_j(G_17_16),.P_i_j(P_17_16));
BlackBlock black_block_19_18(.G_i_k(G_19_19),.P_i_k(P_19_19),.G_km1_j(G_18_18),.P_km1_j(P_18_18),.G_i_j(G_19_18),.P_i_j(P_19_18));
BlackBlock black_block_21_20(.G_i_k(G_21_21),.P_i_k(P_21_21),.G_km1_j(G_20_20),.P_km1_j(P_20_20),.G_i_j(G_21_20),.P_i_j(P_21_20));
BlackBlock black_block_23_22(.G_i_k(G_23_23),.P_i_k(P_23_23),.G_km1_j(G_22_22),.P_km1_j(P_22_22),.G_i_j(G_23_22),.P_i_j(P_23_22));
BlackBlock black_block_25_24(.G_i_k(G_25_25),.P_i_k(P_25_25),.G_km1_j(G_24_24),.P_km1_j(P_24_24),.G_i_j(G_25_24),.P_i_j(P_25_24));
BlackBlock black_block_27_26(.G_i_k(G_27_27),.P_i_k(P_27_27),.G_km1_j(G_26_26),.P_km1_j(P_26_26),.G_i_j(G_27_26),.P_i_j(P_27_26));
BlackBlock black_block_29_28(.G_i_k(G_29_29),.P_i_k(P_29_29),.G_km1_j(G_28_28),.P_km1_j(P_28_28),.G_i_j(G_29_28),.P_i_j(P_29_28));
BlackBlock black_block_31_30(.G_i_k(G_31_31),.P_i_k(P_31_31),.G_km1_j(G_30_30),.P_km1_j(P_30_30),.G_i_j(G_31_30),.P_i_j(P_31_30));
GrayBlock gray_block_3_0(.G_i_k(G_3_2),.P_i_k(P_3_2),.G_km1_j(G_1_0),.G_i_j(G_3_0));
BlackBlock black_block_7_4(.G_i_k(G_7_6),.P_i_k(P_7_6),.G_km1_j(G_5_4),.P_km1_j(P_5_4),.G_i_j(G_7_4),.P_i_j(P_7_4));
BlackBlock black_block_11_8(.G_i_k(G_11_10),.P_i_k(P_11_10),.G_km1_j(G_9_8),.P_km1_j(P_9_8),.G_i_j(G_11_8),.P_i_j(P_11_8));
BlackBlock black_block_15_12(.G_i_k(G_15_14),.P_i_k(P_15_14),.G_km1_j(G_13_12),.P_km1_j(P_13_12),.G_i_j(G_15_12),.P_i_j(P_15_12));
BlackBlock black_block_19_16(.G_i_k(G_19_18),.P_i_k(P_19_18),.G_km1_j(G_17_16),.P_km1_j(P_17_16),.G_i_j(G_19_16),.P_i_j(P_19_16));
BlackBlock black_block_23_20(.G_i_k(G_23_22),.P_i_k(P_23_22),.G_km1_j(G_21_20),.P_km1_j(P_21_20),.G_i_j(G_23_20),.P_i_j(P_23_20));
BlackBlock black_block_27_24(.G_i_k(G_27_26),.P_i_k(P_27_26),.G_km1_j(G_25_24),.P_km1_j(P_25_24),.G_i_j(G_27_24),.P_i_j(P_27_24));
BlackBlock black_block_31_28(.G_i_k(G_31_30),.P_i_k(P_31_30),.G_km1_j(G_29_28),.P_km1_j(P_29_28),.G_i_j(G_31_28),.P_i_j(P_31_28));
GrayBlock gray_block_7_0(.G_i_k(G_7_4),.P_i_k(P_7_4),.G_km1_j(G_3_0),.G_i_j(G_7_0));
BlackBlock black_block_15_8(.G_i_k(G_15_12),.P_i_k(P_15_12),.G_km1_j(G_11_8),.P_km1_j(P_11_8),.G_i_j(G_15_8),.P_i_j(P_15_8));
BlackBlock black_block_23_16(.G_i_k(G_23_20),.P_i_k(P_23_20),.G_km1_j(G_19_16),.P_km1_j(P_19_16),.G_i_j(G_23_16),.P_i_j(P_23_16));
BlackBlock black_block_31_24(.G_i_k(G_31_28),.P_i_k(P_31_28),.G_km1_j(G_27_24),.P_km1_j(P_27_24),.G_i_j(G_31_24),.P_i_j(P_31_24));
GrayBlock gray_block_15_0(.G_i_k(G_15_8),.P_i_k(P_15_8),.G_km1_j(G_7_0),.G_i_j(G_15_0));
BlackBlock black_block_31_16(.G_i_k(G_31_24),.P_i_k(P_31_24),.G_km1_j(G_23_16),.P_km1_j(P_23_16),.G_i_j(G_31_16),.P_i_j(P_31_16));
GrayBlock gray_block_31_0(.G_i_k(G_31_16),.P_i_k(P_31_16),.G_km1_j(G_15_0),.G_i_j(G_31_0));
GrayBlock gray_block_23_15(.G_i_k(G_23_16),.P_i_k(P_23_16),.G_km1_j(G_15_0),.G_i_j(G_23_0));
GrayBlock gray_block_11_7(.G_i_k(G_11_8),.P_i_k(P_11_8),.G_km1_j(G_7_0),.G_i_j(G_11_0));
GrayBlock gray_block_19_15(.G_i_k(G_19_16),.P_i_k(P_19_16),.G_km1_j(G_15_0),.G_i_j(G_19_0));
GrayBlock gray_block_27_23(.G_i_k(G_27_24),.P_i_k(P_27_24),.G_km1_j(G_23_0),.G_i_j(G_27_0));
GrayBlock gray_block_5_3(.G_i_k(G_5_4),.P_i_k(P_5_4),.G_km1_j(G_3_0),.G_i_j(G_5_0));
GrayBlock gray_block_9_7(.G_i_k(G_9_8),.P_i_k(P_9_8),.G_km1_j(G_7_0),.G_i_j(G_9_0));
GrayBlock gray_block_13_11(.G_i_k(G_13_12),.P_i_k(P_13_12),.G_km1_j(G_11_0),.G_i_j(G_13_0));
GrayBlock gray_block_17_15(.G_i_k(G_17_16),.P_i_k(P_17_16),.G_km1_j(G_15_0),.G_i_j(G_17_0));
GrayBlock gray_block_21_19(.G_i_k(G_21_20),.P_i_k(P_21_20),.G_km1_j(G_19_0),.G_i_j(G_21_0));
GrayBlock gray_block_25_23(.G_i_k(G_25_24),.P_i_k(P_25_24),.G_km1_j(G_23_0),.G_i_j(G_25_0));
GrayBlock gray_block_29_27(.G_i_k(G_29_28),.P_i_k(P_29_28),.G_km1_j(G_27_0),.G_i_j(G_29_0));
GrayBlock gray_block_2_1(.G_i_k(G_2_2),.P_i_k(P_2_2),.G_km1_j(G_1_0),.G_i_j(G_2_0));
GrayBlock gray_block_4_3(.G_i_k(G_4_4),.P_i_k(P_4_4),.G_km1_j(G_3_0),.G_i_j(G_4_0));
GrayBlock gray_block_6_5(.G_i_k(G_6_6),.P_i_k(P_6_6),.G_km1_j(G_5_0),.G_i_j(G_6_0));
GrayBlock gray_block_8_7(.G_i_k(G_8_8),.P_i_k(P_8_8),.G_km1_j(G_7_0),.G_i_j(G_8_0));
GrayBlock gray_block_10_9(.G_i_k(G_10_10),.P_i_k(P_10_10),.G_km1_j(G_9_0),.G_i_j(G_10_0));
GrayBlock gray_block_12_11(.G_i_k(G_12_12),.P_i_k(P_12_12),.G_km1_j(G_11_0),.G_i_j(G_12_0));
GrayBlock gray_block_14_13(.G_i_k(G_14_14),.P_i_k(P_14_14),.G_km1_j(G_13_0),.G_i_j(G_14_0));
GrayBlock gray_block_16_15(.G_i_k(G_16_16),.P_i_k(P_16_16),.G_km1_j(G_15_0),.G_i_j(G_16_0));
GrayBlock gray_block_18_17(.G_i_k(G_18_18),.P_i_k(P_18_18),.G_km1_j(G_17_0),.G_i_j(G_18_0));
GrayBlock gray_block_20_19(.G_i_k(G_20_20),.P_i_k(P_20_20),.G_km1_j(G_19_0),.G_i_j(G_20_0));
GrayBlock gray_block_22_21(.G_i_k(G_22_22),.P_i_k(P_22_22),.G_km1_j(G_21_0),.G_i_j(G_22_0));
GrayBlock gray_block_24_23(.G_i_k(G_24_24),.P_i_k(P_24_24),.G_km1_j(G_23_0),.G_i_j(G_24_0));
GrayBlock gray_block_26_25(.G_i_k(G_26_26),.P_i_k(P_26_26),.G_km1_j(G_25_0),.G_i_j(G_26_0));
GrayBlock gray_block_28_27(.G_i_k(G_28_28),.P_i_k(P_28_28),.G_km1_j(G_27_0),.G_i_j(G_28_0));
GrayBlock gray_block_30_29(.G_i_k(G_30_30),.P_i_k(P_30_30),.G_km1_j(G_29_0),.G_i_j(G_30_0));
GrayBlock gray_block_32_31(.G_i_k(G_32_32),.P_i_k(P_32_32),.G_km1_j(G_31_0),.G_i_j(G_32_0));
assign _P_0_0 = P_0_0 ;
assign _G_0_0 = G_0_0 ;
endmodule
