module BrentKungAdder ( A_1,B_1,A_2,B_2,A_3,B_3,A_4,B_4,A_5,B_5,A_6,B_6,A_7,B_7,A_8,B_8,C_0,S_1,S_2,S_3,S_4,S_5,S_6,S_7,S_8,C_out );
input A_1;
input B_1;
input A_2;
input B_2;
input A_3;
input B_3;
input A_4;
input B_4;
input A_5;
input B_5;
input A_6;
input B_6;
input A_7;
input B_7;
input A_8;
input B_8;
input C_0;
output S_1;
output S_2;
output S_3;
output S_4;
output S_5;
output S_6;
output S_7;
output S_8;
output C_out;
wire P_0;
wire G_0;
wire P_1;
wire G_1;
wire P_2;
wire G_2;
wire P_3;
wire G_3;
wire P_4;
wire G_4;
wire P_5;
wire G_5;
wire P_6;
wire G_6;
wire P_7;
wire G_7;
wire P_8;
wire G_8;
wire P_0_0;
wire G_0_0;
wire P_1_0;
wire G_1_0;
wire P_2_0;
wire G_2_0;
wire P_3_0;
wire G_3_0;
wire P_4_0;
wire G_4_0;
wire P_5_0;
wire G_5_0;
wire P_6_0;
wire G_6_0;
wire P_7_0;
wire G_7_0;
wire P_8_0;
wire G_8_0;
BitwisePGLogic _BitwisePGLogic(.C_0(C_0),.A_1(A_1),.B_1(B_1),.A_2(A_2),.B_2(B_2),.A_3(A_3),.B_3(B_3),.A_4(A_4),.B_4(B_4),.A_5(A_5),.B_5(B_5),.A_6(A_6),.B_6(B_6),.A_7(A_7),.B_7(B_7),.A_8(A_8),.B_8(B_8),.P_0(P_0),.G_0(G_0),.P_1(P_1),.G_1(G_1),.P_2(P_2),.G_2(G_2),.P_3(P_3),.G_3(G_3),.P_4(P_4),.G_4(G_4),.P_5(P_5),.G_5(G_5),.P_6(P_6),.G_6(G_6),.P_7(P_7),.G_7(G_7),.P_8(P_8),.G_8(G_8));
GroupPGLogic _GroupPGLogic(.P_0_0(P_0),.G_0_0(G_0),.P_1_1(P_1),.G_1_1(G_1),.P_2_2(P_2),.G_2_2(G_2),.P_3_3(P_3),.G_3_3(G_3),.P_4_4(P_4),.G_4_4(G_4),.P_5_5(P_5),.G_5_5(G_5),.P_6_6(P_6),.G_6_6(G_6),.P_7_7(P_7),.G_7_7(G_7),.P_8_8(P_8),.G_8_8(G_8),._P_0_0(P_0_0),._G_0_0(G_0_0),.P_1_0(P_1_0),.G_1_0(G_1_0),.P_2_0(P_2_0),.G_2_0(G_2_0),.P_3_0(P_3_0),.G_3_0(G_3_0),.P_4_0(P_4_0),.G_4_0(G_4_0),.P_5_0(P_5_0),.G_5_0(G_5_0),.P_6_0(P_6_0),.G_6_0(G_6_0),.P_7_0(P_7_0),.G_7_0(G_7_0),.P_8_0(P_8_0),.G_8_0(G_8_0));
SumLogic _SumLogic(.P_0(P_0),.G_0_0(G_0_0),.P_1(P_1),.G_1_0(G_1_0),.P_2(P_2),.G_2_0(G_2_0),.P_3(P_3),.G_3_0(G_3_0),.P_4(P_4),.G_4_0(G_4_0),.P_5(P_5),.G_5_0(G_5_0),.P_6(P_6),.G_6_0(G_6_0),.P_7(P_7),.G_7_0(G_7_0),.P_8(P_8),.G_8_0(G_8_0),.S_1(S_1),.S_2(S_2),.S_3(S_3),.S_4(S_4),.S_5(S_5),.S_6(S_6),.S_7(S_7),.S_8(S_8),.C_out(C_out));
endmodule
