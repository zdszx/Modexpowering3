module BitwisePGLogic ( A_1,B_1,A_2,B_2,A_3,B_3,A_4,B_4,A_5,B_5,A_6,B_6,A_7,B_7,A_8,B_8,A_9,B_9,A_10,B_10,A_11,B_11,A_12,B_12,A_13,B_13,A_14,B_14,A_15,B_15,A_16,B_16,A_17,B_17,A_18,B_18,A_19,B_19,A_20,B_20,A_21,B_21,A_22,B_22,A_23,B_23,A_24,B_24,A_25,B_25,A_26,B_26,A_27,B_27,A_28,B_28,A_29,B_29,A_30,B_30,A_31,B_31,A_32,B_32,C_0,P_0,G_0,P_1,G_1,P_2,G_2,P_3,G_3,P_4,G_4,P_5,G_5,P_6,G_6,P_7,G_7,P_8,G_8,P_9,G_9,P_10,G_10,P_11,G_11,P_12,G_12,P_13,G_13,P_14,G_14,P_15,G_15,P_16,G_16,P_17,G_17,P_18,G_18,P_19,G_19,P_20,G_20,P_21,G_21,P_22,G_22,P_23,G_23,P_24,G_24,P_25,G_25,P_26,G_26,P_27,G_27,P_28,G_28,P_29,G_29,P_30,G_30,P_31,G_31,P_32,G_32 );
input A_1;
input B_1;
input A_2;
input B_2;
input A_3;
input B_3;
input A_4;
input B_4;
input A_5;
input B_5;
input A_6;
input B_6;
input A_7;
input B_7;
input A_8;
input B_8;
input A_9;
input B_9;
input A_10;
input B_10;
input A_11;
input B_11;
input A_12;
input B_12;
input A_13;
input B_13;
input A_14;
input B_14;
input A_15;
input B_15;
input A_16;
input B_16;
input A_17;
input B_17;
input A_18;
input B_18;
input A_19;
input B_19;
input A_20;
input B_20;
input A_21;
input B_21;
input A_22;
input B_22;
input A_23;
input B_23;
input A_24;
input B_24;
input A_25;
input B_25;
input A_26;
input B_26;
input A_27;
input B_27;
input A_28;
input B_28;
input A_29;
input B_29;
input A_30;
input B_30;
input A_31;
input B_31;
input A_32;
input B_32;
input C_0;
output P_0;
output G_0;
output P_1;
output G_1;
output P_2;
output G_2;
output P_3;
output G_3;
output P_4;
output G_4;
output P_5;
output G_5;
output P_6;
output G_6;
output P_7;
output G_7;
output P_8;
output G_8;
output P_9;
output G_9;
output P_10;
output G_10;
output P_11;
output G_11;
output P_12;
output G_12;
output P_13;
output G_13;
output P_14;
output G_14;
output P_15;
output G_15;
output P_16;
output G_16;
output P_17;
output G_17;
output P_18;
output G_18;
output P_19;
output G_19;
output P_20;
output G_20;
output P_21;
output G_21;
output P_22;
output G_22;
output P_23;
output G_23;
output P_24;
output G_24;
output P_25;
output G_25;
output P_26;
output G_26;
output P_27;
output G_27;
output P_28;
output G_28;
output P_29;
output G_29;
output P_30;
output G_30;
output P_31;
output G_31;
output P_32;
output G_32;
// Bit 0
assign P_0 = 0 ;
assign G_0 = C_0 ;
// Bit 1
PG PG_Bit_1(.A_i(A_1),.B_i(B_1),.P_i(P_1),.G_i(G_1));
// Bit 2
PG PG_Bit_2(.A_i(A_2),.B_i(B_2),.P_i(P_2),.G_i(G_2));
// Bit 3
PG PG_Bit_3(.A_i(A_3),.B_i(B_3),.P_i(P_3),.G_i(G_3));
// Bit 4
PG PG_Bit_4(.A_i(A_4),.B_i(B_4),.P_i(P_4),.G_i(G_4));
// Bit 5
PG PG_Bit_5(.A_i(A_5),.B_i(B_5),.P_i(P_5),.G_i(G_5));
// Bit 6
PG PG_Bit_6(.A_i(A_6),.B_i(B_6),.P_i(P_6),.G_i(G_6));
// Bit 7
PG PG_Bit_7(.A_i(A_7),.B_i(B_7),.P_i(P_7),.G_i(G_7));
// Bit 8
PG PG_Bit_8(.A_i(A_8),.B_i(B_8),.P_i(P_8),.G_i(G_8));
// Bit 9
PG PG_Bit_9(.A_i(A_9),.B_i(B_9),.P_i(P_9),.G_i(G_9));
// Bit 10
PG PG_Bit_10(.A_i(A_10),.B_i(B_10),.P_i(P_10),.G_i(G_10));
// Bit 11
PG PG_Bit_11(.A_i(A_11),.B_i(B_11),.P_i(P_11),.G_i(G_11));
// Bit 12
PG PG_Bit_12(.A_i(A_12),.B_i(B_12),.P_i(P_12),.G_i(G_12));
// Bit 13
PG PG_Bit_13(.A_i(A_13),.B_i(B_13),.P_i(P_13),.G_i(G_13));
// Bit 14
PG PG_Bit_14(.A_i(A_14),.B_i(B_14),.P_i(P_14),.G_i(G_14));
// Bit 15
PG PG_Bit_15(.A_i(A_15),.B_i(B_15),.P_i(P_15),.G_i(G_15));
// Bit 16
PG PG_Bit_16(.A_i(A_16),.B_i(B_16),.P_i(P_16),.G_i(G_16));
// Bit 17
PG PG_Bit_17(.A_i(A_17),.B_i(B_17),.P_i(P_17),.G_i(G_17));
// Bit 18
PG PG_Bit_18(.A_i(A_18),.B_i(B_18),.P_i(P_18),.G_i(G_18));
// Bit 19
PG PG_Bit_19(.A_i(A_19),.B_i(B_19),.P_i(P_19),.G_i(G_19));
// Bit 20
PG PG_Bit_20(.A_i(A_20),.B_i(B_20),.P_i(P_20),.G_i(G_20));
// Bit 21
PG PG_Bit_21(.A_i(A_21),.B_i(B_21),.P_i(P_21),.G_i(G_21));
// Bit 22
PG PG_Bit_22(.A_i(A_22),.B_i(B_22),.P_i(P_22),.G_i(G_22));
// Bit 23
PG PG_Bit_23(.A_i(A_23),.B_i(B_23),.P_i(P_23),.G_i(G_23));
// Bit 24
PG PG_Bit_24(.A_i(A_24),.B_i(B_24),.P_i(P_24),.G_i(G_24));
// Bit 25
PG PG_Bit_25(.A_i(A_25),.B_i(B_25),.P_i(P_25),.G_i(G_25));
// Bit 26
PG PG_Bit_26(.A_i(A_26),.B_i(B_26),.P_i(P_26),.G_i(G_26));
// Bit 27
PG PG_Bit_27(.A_i(A_27),.B_i(B_27),.P_i(P_27),.G_i(G_27));
// Bit 28
PG PG_Bit_28(.A_i(A_28),.B_i(B_28),.P_i(P_28),.G_i(G_28));
// Bit 29
PG PG_Bit_29(.A_i(A_29),.B_i(B_29),.P_i(P_29),.G_i(G_29));
// Bit 30
PG PG_Bit_30(.A_i(A_30),.B_i(B_30),.P_i(P_30),.G_i(G_30));
// Bit 31
PG PG_Bit_31(.A_i(A_31),.B_i(B_31),.P_i(P_31),.G_i(G_31));
// Bit 32
PG PG_Bit_32(.A_i(A_32),.B_i(B_32),.P_i(P_32),.G_i(G_32));
endmodule
