module GroupPGLogic ( P_0_0,G_0_0,P_1_1,G_1_1,P_2_2,G_2_2,P_3_3,G_3_3,P_4_4,G_4_4,_P_0_0,_G_0_0,P_1_0,G_1_0,P_2_0,G_2_0,P_3_0,G_3_0,P_4_0,G_4_0 );
input P_0_0;
input G_0_0;
input P_1_1;
input G_1_1;
input P_2_2;
input G_2_2;
input P_3_3;
input G_3_3;
input P_4_4;
input G_4_4;
output _P_0_0;
output _G_0_0;
output P_1_0;
output G_1_0;
output P_2_0;
output G_2_0;
output P_3_0;
output G_3_0;
output P_4_0;
output G_4_0;
wire G_3_2;
wire P_3_2;
GrayBlock gray_block_1_0(.G_i_k(G_1_1),.P_i_k(P_1_1),.G_km1_j(G_0_0),.G_i_j(G_1_0));
BlackBlock black_block_3_2(.G_i_k(G_3_3),.P_i_k(P_3_3),.G_km1_j(G_2_2),.P_km1_j(P_2_2),.G_i_j(G_3_2),.P_i_j(P_3_2));
GrayBlock gray_block_3_0(.G_i_k(G_3_2),.P_i_k(P_3_2),.G_km1_j(G_1_0),.G_i_j(G_3_0));
GrayBlock gray_block_2_1(.G_i_k(G_2_2),.P_i_k(P_2_2),.G_km1_j(G_1_0),.G_i_j(G_2_0));
GrayBlock gray_block_4_3(.G_i_k(G_4_4),.P_i_k(P_4_4),.G_km1_j(G_3_0),.G_i_j(G_4_0));
assign _P_0_0 = P_0_0 ;
assign _G_0_0 = G_0_0 ;
endmodule
