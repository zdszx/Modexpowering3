module SumLogic ( P_0,G_0_0,P_1,G_1_0,P_2,G_2_0,P_3,G_3_0,P_4,G_4_0,P_5,G_5_0,P_6,G_6_0,P_7,G_7_0,P_8,G_8_0,P_9,G_9_0,P_10,G_10_0,P_11,G_11_0,P_12,G_12_0,P_13,G_13_0,P_14,G_14_0,P_15,G_15_0,P_16,G_16_0,P_17,G_17_0,P_18,G_18_0,P_19,G_19_0,P_20,G_20_0,P_21,G_21_0,P_22,G_22_0,P_23,G_23_0,P_24,G_24_0,P_25,G_25_0,P_26,G_26_0,P_27,G_27_0,P_28,G_28_0,P_29,G_29_0,P_30,G_30_0,P_31,G_31_0,P_32,G_32_0,S_1,S_2,S_3,S_4,S_5,S_6,S_7,S_8,S_9,S_10,S_11,S_12,S_13,S_14,S_15,S_16,S_17,S_18,S_19,S_20,S_21,S_22,S_23,S_24,S_25,S_26,S_27,S_28,S_29,S_30,S_31,S_32,C_out );
input P_0;
input G_0_0;
input P_1;
input G_1_0;
input P_2;
input G_2_0;
input P_3;
input G_3_0;
input P_4;
input G_4_0;
input P_5;
input G_5_0;
input P_6;
input G_6_0;
input P_7;
input G_7_0;
input P_8;
input G_8_0;
input P_9;
input G_9_0;
input P_10;
input G_10_0;
input P_11;
input G_11_0;
input P_12;
input G_12_0;
input P_13;
input G_13_0;
input P_14;
input G_14_0;
input P_15;
input G_15_0;
input P_16;
input G_16_0;
input P_17;
input G_17_0;
input P_18;
input G_18_0;
input P_19;
input G_19_0;
input P_20;
input G_20_0;
input P_21;
input G_21_0;
input P_22;
input G_22_0;
input P_23;
input G_23_0;
input P_24;
input G_24_0;
input P_25;
input G_25_0;
input P_26;
input G_26_0;
input P_27;
input G_27_0;
input P_28;
input G_28_0;
input P_29;
input G_29_0;
input P_30;
input G_30_0;
input P_31;
input G_31_0;
input P_32;
input G_32_0;
output S_1;
output S_2;
output S_3;
output S_4;
output S_5;
output S_6;
output S_7;
output S_8;
output S_9;
output S_10;
output S_11;
output S_12;
output S_13;
output S_14;
output S_15;
output S_16;
output S_17;
output S_18;
output S_19;
output S_20;
output S_21;
output S_22;
output S_23;
output S_24;
output S_25;
output S_26;
output S_27;
output S_28;
output S_29;
output S_30;
output S_31;
output S_32;
output C_out;
// Bit 1
assign S_1 = G_0_0 ^ P_1 ;
// Bit 2
assign S_2 = G_1_0 ^ P_2 ;
// Bit 3
assign S_3 = G_2_0 ^ P_3 ;
// Bit 4
assign S_4 = G_3_0 ^ P_4 ;
// Bit 5
assign S_5 = G_4_0 ^ P_5 ;
// Bit 6
assign S_6 = G_5_0 ^ P_6 ;
// Bit 7
assign S_7 = G_6_0 ^ P_7 ;
// Bit 8
assign S_8 = G_7_0 ^ P_8 ;
// Bit 9
assign S_9 = G_8_0 ^ P_9 ;
// Bit 10
assign S_10 = G_9_0 ^ P_10 ;
// Bit 11
assign S_11 = G_10_0 ^ P_11 ;
// Bit 12
assign S_12 = G_11_0 ^ P_12 ;
// Bit 13
assign S_13 = G_12_0 ^ P_13 ;
// Bit 14
assign S_14 = G_13_0 ^ P_14 ;
// Bit 15
assign S_15 = G_14_0 ^ P_15 ;
// Bit 16
assign S_16 = G_15_0 ^ P_16 ;
// Bit 17
assign S_17 = G_16_0 ^ P_17 ;
// Bit 18
assign S_18 = G_17_0 ^ P_18 ;
// Bit 19
assign S_19 = G_18_0 ^ P_19 ;
// Bit 20
assign S_20 = G_19_0 ^ P_20 ;
// Bit 21
assign S_21 = G_20_0 ^ P_21 ;
// Bit 22
assign S_22 = G_21_0 ^ P_22 ;
// Bit 23
assign S_23 = G_22_0 ^ P_23 ;
// Bit 24
assign S_24 = G_23_0 ^ P_24 ;
// Bit 25
assign S_25 = G_24_0 ^ P_25 ;
// Bit 26
assign S_26 = G_25_0 ^ P_26 ;
// Bit 27
assign S_27 = G_26_0 ^ P_27 ;
// Bit 28
assign S_28 = G_27_0 ^ P_28 ;
// Bit 29
assign S_29 = G_28_0 ^ P_29 ;
// Bit 30
assign S_30 = G_29_0 ^ P_30 ;
// Bit 31
assign S_31 = G_30_0 ^ P_31 ;
// Bit 32
assign S_32 = G_31_0 ^ P_32 ;
// Carry Out
assign C_out = G_32_0 ;
endmodule
