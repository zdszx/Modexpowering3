module SumLogic ( P_0,G_0_0,P_1,G_1_0,P_2,G_2_0,P_3,G_3_0,P_4,G_4_0,P_5,G_5_0,P_6,G_6_0,P_7,G_7_0,P_8,G_8_0,P_9,G_9_0,P_10,G_10_0,P_11,G_11_0,P_12,G_12_0,P_13,G_13_0,P_14,G_14_0,P_15,G_15_0,P_16,G_16_0,P_17,G_17_0,P_18,G_18_0,P_19,G_19_0,P_20,G_20_0,P_21,G_21_0,P_22,G_22_0,P_23,G_23_0,P_24,G_24_0,P_25,G_25_0,P_26,G_26_0,P_27,G_27_0,P_28,G_28_0,P_29,G_29_0,P_30,G_30_0,P_31,G_31_0,P_32,G_32_0,P_33,G_33_0,P_34,G_34_0,P_35,G_35_0,P_36,G_36_0,P_37,G_37_0,P_38,G_38_0,P_39,G_39_0,P_40,G_40_0,P_41,G_41_0,P_42,G_42_0,P_43,G_43_0,P_44,G_44_0,P_45,G_45_0,P_46,G_46_0,P_47,G_47_0,P_48,G_48_0,P_49,G_49_0,P_50,G_50_0,P_51,G_51_0,P_52,G_52_0,P_53,G_53_0,P_54,G_54_0,P_55,G_55_0,P_56,G_56_0,P_57,G_57_0,P_58,G_58_0,P_59,G_59_0,P_60,G_60_0,P_61,G_61_0,P_62,G_62_0,P_63,G_63_0,P_64,G_64_0,S_1,S_2,S_3,S_4,S_5,S_6,S_7,S_8,S_9,S_10,S_11,S_12,S_13,S_14,S_15,S_16,S_17,S_18,S_19,S_20,S_21,S_22,S_23,S_24,S_25,S_26,S_27,S_28,S_29,S_30,S_31,S_32,S_33,S_34,S_35,S_36,S_37,S_38,S_39,S_40,S_41,S_42,S_43,S_44,S_45,S_46,S_47,S_48,S_49,S_50,S_51,S_52,S_53,S_54,S_55,S_56,S_57,S_58,S_59,S_60,S_61,S_62,S_63,S_64,C_out );
input P_0;
input G_0_0;
input P_1;
input G_1_0;
input P_2;
input G_2_0;
input P_3;
input G_3_0;
input P_4;
input G_4_0;
input P_5;
input G_5_0;
input P_6;
input G_6_0;
input P_7;
input G_7_0;
input P_8;
input G_8_0;
input P_9;
input G_9_0;
input P_10;
input G_10_0;
input P_11;
input G_11_0;
input P_12;
input G_12_0;
input P_13;
input G_13_0;
input P_14;
input G_14_0;
input P_15;
input G_15_0;
input P_16;
input G_16_0;
input P_17;
input G_17_0;
input P_18;
input G_18_0;
input P_19;
input G_19_0;
input P_20;
input G_20_0;
input P_21;
input G_21_0;
input P_22;
input G_22_0;
input P_23;
input G_23_0;
input P_24;
input G_24_0;
input P_25;
input G_25_0;
input P_26;
input G_26_0;
input P_27;
input G_27_0;
input P_28;
input G_28_0;
input P_29;
input G_29_0;
input P_30;
input G_30_0;
input P_31;
input G_31_0;
input P_32;
input G_32_0;
input P_33;
input G_33_0;
input P_34;
input G_34_0;
input P_35;
input G_35_0;
input P_36;
input G_36_0;
input P_37;
input G_37_0;
input P_38;
input G_38_0;
input P_39;
input G_39_0;
input P_40;
input G_40_0;
input P_41;
input G_41_0;
input P_42;
input G_42_0;
input P_43;
input G_43_0;
input P_44;
input G_44_0;
input P_45;
input G_45_0;
input P_46;
input G_46_0;
input P_47;
input G_47_0;
input P_48;
input G_48_0;
input P_49;
input G_49_0;
input P_50;
input G_50_0;
input P_51;
input G_51_0;
input P_52;
input G_52_0;
input P_53;
input G_53_0;
input P_54;
input G_54_0;
input P_55;
input G_55_0;
input P_56;
input G_56_0;
input P_57;
input G_57_0;
input P_58;
input G_58_0;
input P_59;
input G_59_0;
input P_60;
input G_60_0;
input P_61;
input G_61_0;
input P_62;
input G_62_0;
input P_63;
input G_63_0;
input P_64;
input G_64_0;
output S_1;
output S_2;
output S_3;
output S_4;
output S_5;
output S_6;
output S_7;
output S_8;
output S_9;
output S_10;
output S_11;
output S_12;
output S_13;
output S_14;
output S_15;
output S_16;
output S_17;
output S_18;
output S_19;
output S_20;
output S_21;
output S_22;
output S_23;
output S_24;
output S_25;
output S_26;
output S_27;
output S_28;
output S_29;
output S_30;
output S_31;
output S_32;
output S_33;
output S_34;
output S_35;
output S_36;
output S_37;
output S_38;
output S_39;
output S_40;
output S_41;
output S_42;
output S_43;
output S_44;
output S_45;
output S_46;
output S_47;
output S_48;
output S_49;
output S_50;
output S_51;
output S_52;
output S_53;
output S_54;
output S_55;
output S_56;
output S_57;
output S_58;
output S_59;
output S_60;
output S_61;
output S_62;
output S_63;
output S_64;
output C_out;
// Bit 1
assign S_1 = G_0_0 ^ P_1 ;
// Bit 2
assign S_2 = G_1_0 ^ P_2 ;
// Bit 3
assign S_3 = G_2_0 ^ P_3 ;
// Bit 4
assign S_4 = G_3_0 ^ P_4 ;
// Bit 5
assign S_5 = G_4_0 ^ P_5 ;
// Bit 6
assign S_6 = G_5_0 ^ P_6 ;
// Bit 7
assign S_7 = G_6_0 ^ P_7 ;
// Bit 8
assign S_8 = G_7_0 ^ P_8 ;
// Bit 9
assign S_9 = G_8_0 ^ P_9 ;
// Bit 10
assign S_10 = G_9_0 ^ P_10 ;
// Bit 11
assign S_11 = G_10_0 ^ P_11 ;
// Bit 12
assign S_12 = G_11_0 ^ P_12 ;
// Bit 13
assign S_13 = G_12_0 ^ P_13 ;
// Bit 14
assign S_14 = G_13_0 ^ P_14 ;
// Bit 15
assign S_15 = G_14_0 ^ P_15 ;
// Bit 16
assign S_16 = G_15_0 ^ P_16 ;
// Bit 17
assign S_17 = G_16_0 ^ P_17 ;
// Bit 18
assign S_18 = G_17_0 ^ P_18 ;
// Bit 19
assign S_19 = G_18_0 ^ P_19 ;
// Bit 20
assign S_20 = G_19_0 ^ P_20 ;
// Bit 21
assign S_21 = G_20_0 ^ P_21 ;
// Bit 22
assign S_22 = G_21_0 ^ P_22 ;
// Bit 23
assign S_23 = G_22_0 ^ P_23 ;
// Bit 24
assign S_24 = G_23_0 ^ P_24 ;
// Bit 25
assign S_25 = G_24_0 ^ P_25 ;
// Bit 26
assign S_26 = G_25_0 ^ P_26 ;
// Bit 27
assign S_27 = G_26_0 ^ P_27 ;
// Bit 28
assign S_28 = G_27_0 ^ P_28 ;
// Bit 29
assign S_29 = G_28_0 ^ P_29 ;
// Bit 30
assign S_30 = G_29_0 ^ P_30 ;
// Bit 31
assign S_31 = G_30_0 ^ P_31 ;
// Bit 32
assign S_32 = G_31_0 ^ P_32 ;
// Bit 33
assign S_33 = G_32_0 ^ P_33 ;
// Bit 34
assign S_34 = G_33_0 ^ P_34 ;
// Bit 35
assign S_35 = G_34_0 ^ P_35 ;
// Bit 36
assign S_36 = G_35_0 ^ P_36 ;
// Bit 37
assign S_37 = G_36_0 ^ P_37 ;
// Bit 38
assign S_38 = G_37_0 ^ P_38 ;
// Bit 39
assign S_39 = G_38_0 ^ P_39 ;
// Bit 40
assign S_40 = G_39_0 ^ P_40 ;
// Bit 41
assign S_41 = G_40_0 ^ P_41 ;
// Bit 42
assign S_42 = G_41_0 ^ P_42 ;
// Bit 43
assign S_43 = G_42_0 ^ P_43 ;
// Bit 44
assign S_44 = G_43_0 ^ P_44 ;
// Bit 45
assign S_45 = G_44_0 ^ P_45 ;
// Bit 46
assign S_46 = G_45_0 ^ P_46 ;
// Bit 47
assign S_47 = G_46_0 ^ P_47 ;
// Bit 48
assign S_48 = G_47_0 ^ P_48 ;
// Bit 49
assign S_49 = G_48_0 ^ P_49 ;
// Bit 50
assign S_50 = G_49_0 ^ P_50 ;
// Bit 51
assign S_51 = G_50_0 ^ P_51 ;
// Bit 52
assign S_52 = G_51_0 ^ P_52 ;
// Bit 53
assign S_53 = G_52_0 ^ P_53 ;
// Bit 54
assign S_54 = G_53_0 ^ P_54 ;
// Bit 55
assign S_55 = G_54_0 ^ P_55 ;
// Bit 56
assign S_56 = G_55_0 ^ P_56 ;
// Bit 57
assign S_57 = G_56_0 ^ P_57 ;
// Bit 58
assign S_58 = G_57_0 ^ P_58 ;
// Bit 59
assign S_59 = G_58_0 ^ P_59 ;
// Bit 60
assign S_60 = G_59_0 ^ P_60 ;
// Bit 61
assign S_61 = G_60_0 ^ P_61 ;
// Bit 62
assign S_62 = G_61_0 ^ P_62 ;
// Bit 63
assign S_63 = G_62_0 ^ P_63 ;
// Bit 64
assign S_64 = G_63_0 ^ P_64 ;
// Carry Out
assign C_out = G_64_0 ;
endmodule
