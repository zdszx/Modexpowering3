module BrentKungAdder ( A_1,B_1,A_2,B_2,A_3,B_3,A_4,B_4,A_5,B_5,A_6,B_6,A_7,B_7,A_8,B_8,A_9,B_9,A_10,B_10,A_11,B_11,A_12,B_12,A_13,B_13,A_14,B_14,A_15,B_15,A_16,B_16,A_17,B_17,A_18,B_18,A_19,B_19,A_20,B_20,A_21,B_21,A_22,B_22,A_23,B_23,A_24,B_24,A_25,B_25,A_26,B_26,A_27,B_27,A_28,B_28,A_29,B_29,A_30,B_30,A_31,B_31,A_32,B_32,C_0,S_1,S_2,S_3,S_4,S_5,S_6,S_7,S_8,S_9,S_10,S_11,S_12,S_13,S_14,S_15,S_16,S_17,S_18,S_19,S_20,S_21,S_22,S_23,S_24,S_25,S_26,S_27,S_28,S_29,S_30,S_31,S_32,C_out );
input A_1;
input B_1;
input A_2;
input B_2;
input A_3;
input B_3;
input A_4;
input B_4;
input A_5;
input B_5;
input A_6;
input B_6;
input A_7;
input B_7;
input A_8;
input B_8;
input A_9;
input B_9;
input A_10;
input B_10;
input A_11;
input B_11;
input A_12;
input B_12;
input A_13;
input B_13;
input A_14;
input B_14;
input A_15;
input B_15;
input A_16;
input B_16;
input A_17;
input B_17;
input A_18;
input B_18;
input A_19;
input B_19;
input A_20;
input B_20;
input A_21;
input B_21;
input A_22;
input B_22;
input A_23;
input B_23;
input A_24;
input B_24;
input A_25;
input B_25;
input A_26;
input B_26;
input A_27;
input B_27;
input A_28;
input B_28;
input A_29;
input B_29;
input A_30;
input B_30;
input A_31;
input B_31;
input A_32;
input B_32;
input C_0;
output S_1;
output S_2;
output S_3;
output S_4;
output S_5;
output S_6;
output S_7;
output S_8;
output S_9;
output S_10;
output S_11;
output S_12;
output S_13;
output S_14;
output S_15;
output S_16;
output S_17;
output S_18;
output S_19;
output S_20;
output S_21;
output S_22;
output S_23;
output S_24;
output S_25;
output S_26;
output S_27;
output S_28;
output S_29;
output S_30;
output S_31;
output S_32;
output C_out;
wire P_0;
wire G_0;
wire P_1;
wire G_1;
wire P_2;
wire G_2;
wire P_3;
wire G_3;
wire P_4;
wire G_4;
wire P_5;
wire G_5;
wire P_6;
wire G_6;
wire P_7;
wire G_7;
wire P_8;
wire G_8;
wire P_9;
wire G_9;
wire P_10;
wire G_10;
wire P_11;
wire G_11;
wire P_12;
wire G_12;
wire P_13;
wire G_13;
wire P_14;
wire G_14;
wire P_15;
wire G_15;
wire P_16;
wire G_16;
wire P_17;
wire G_17;
wire P_18;
wire G_18;
wire P_19;
wire G_19;
wire P_20;
wire G_20;
wire P_21;
wire G_21;
wire P_22;
wire G_22;
wire P_23;
wire G_23;
wire P_24;
wire G_24;
wire P_25;
wire G_25;
wire P_26;
wire G_26;
wire P_27;
wire G_27;
wire P_28;
wire G_28;
wire P_29;
wire G_29;
wire P_30;
wire G_30;
wire P_31;
wire G_31;
wire P_32;
wire G_32;
wire P_0_0;
wire G_0_0;
wire P_1_0;
wire G_1_0;
wire P_2_0;
wire G_2_0;
wire P_3_0;
wire G_3_0;
wire P_4_0;
wire G_4_0;
wire P_5_0;
wire G_5_0;
wire P_6_0;
wire G_6_0;
wire P_7_0;
wire G_7_0;
wire P_8_0;
wire G_8_0;
wire P_9_0;
wire G_9_0;
wire P_10_0;
wire G_10_0;
wire P_11_0;
wire G_11_0;
wire P_12_0;
wire G_12_0;
wire P_13_0;
wire G_13_0;
wire P_14_0;
wire G_14_0;
wire P_15_0;
wire G_15_0;
wire P_16_0;
wire G_16_0;
wire P_17_0;
wire G_17_0;
wire P_18_0;
wire G_18_0;
wire P_19_0;
wire G_19_0;
wire P_20_0;
wire G_20_0;
wire P_21_0;
wire G_21_0;
wire P_22_0;
wire G_22_0;
wire P_23_0;
wire G_23_0;
wire P_24_0;
wire G_24_0;
wire P_25_0;
wire G_25_0;
wire P_26_0;
wire G_26_0;
wire P_27_0;
wire G_27_0;
wire P_28_0;
wire G_28_0;
wire P_29_0;
wire G_29_0;
wire P_30_0;
wire G_30_0;
wire P_31_0;
wire G_31_0;
wire P_32_0;
wire G_32_0;
BitwisePGLogic _BitwisePGLogic(.C_0(C_0),.A_1(A_1),.B_1(B_1),.A_2(A_2),.B_2(B_2),.A_3(A_3),.B_3(B_3),.A_4(A_4),.B_4(B_4),.A_5(A_5),.B_5(B_5),.A_6(A_6),.B_6(B_6),.A_7(A_7),.B_7(B_7),.A_8(A_8),.B_8(B_8),.A_9(A_9),.B_9(B_9),.A_10(A_10),.B_10(B_10),.A_11(A_11),.B_11(B_11),.A_12(A_12),.B_12(B_12),.A_13(A_13),.B_13(B_13),.A_14(A_14),.B_14(B_14),.A_15(A_15),.B_15(B_15),.A_16(A_16),.B_16(B_16),.A_17(A_17),.B_17(B_17),.A_18(A_18),.B_18(B_18),.A_19(A_19),.B_19(B_19),.A_20(A_20),.B_20(B_20),.A_21(A_21),.B_21(B_21),.A_22(A_22),.B_22(B_22),.A_23(A_23),.B_23(B_23),.A_24(A_24),.B_24(B_24),.A_25(A_25),.B_25(B_25),.A_26(A_26),.B_26(B_26),.A_27(A_27),.B_27(B_27),.A_28(A_28),.B_28(B_28),.A_29(A_29),.B_29(B_29),.A_30(A_30),.B_30(B_30),.A_31(A_31),.B_31(B_31),.A_32(A_32),.B_32(B_32),.P_0(P_0),.G_0(G_0),.P_1(P_1),.G_1(G_1),.P_2(P_2),.G_2(G_2),.P_3(P_3),.G_3(G_3),.P_4(P_4),.G_4(G_4),.P_5(P_5),.G_5(G_5),.P_6(P_6),.G_6(G_6),.P_7(P_7),.G_7(G_7),.P_8(P_8),.G_8(G_8),.P_9(P_9),.G_9(G_9),.P_10(P_10),.G_10(G_10),.P_11(P_11),.G_11(G_11),.P_12(P_12),.G_12(G_12),.P_13(P_13),.G_13(G_13),.P_14(P_14),.G_14(G_14),.P_15(P_15),.G_15(G_15),.P_16(P_16),.G_16(G_16),.P_17(P_17),.G_17(G_17),.P_18(P_18),.G_18(G_18),.P_19(P_19),.G_19(G_19),.P_20(P_20),.G_20(G_20),.P_21(P_21),.G_21(G_21),.P_22(P_22),.G_22(G_22),.P_23(P_23),.G_23(G_23),.P_24(P_24),.G_24(G_24),.P_25(P_25),.G_25(G_25),.P_26(P_26),.G_26(G_26),.P_27(P_27),.G_27(G_27),.P_28(P_28),.G_28(G_28),.P_29(P_29),.G_29(G_29),.P_30(P_30),.G_30(G_30),.P_31(P_31),.G_31(G_31),.P_32(P_32),.G_32(G_32));
GroupPGLogic _GroupPGLogic(.P_0_0(P_0),.G_0_0(G_0),.P_1_1(P_1),.G_1_1(G_1),.P_2_2(P_2),.G_2_2(G_2),.P_3_3(P_3),.G_3_3(G_3),.P_4_4(P_4),.G_4_4(G_4),.P_5_5(P_5),.G_5_5(G_5),.P_6_6(P_6),.G_6_6(G_6),.P_7_7(P_7),.G_7_7(G_7),.P_8_8(P_8),.G_8_8(G_8),.P_9_9(P_9),.G_9_9(G_9),.P_10_10(P_10),.G_10_10(G_10),.P_11_11(P_11),.G_11_11(G_11),.P_12_12(P_12),.G_12_12(G_12),.P_13_13(P_13),.G_13_13(G_13),.P_14_14(P_14),.G_14_14(G_14),.P_15_15(P_15),.G_15_15(G_15),.P_16_16(P_16),.G_16_16(G_16),.P_17_17(P_17),.G_17_17(G_17),.P_18_18(P_18),.G_18_18(G_18),.P_19_19(P_19),.G_19_19(G_19),.P_20_20(P_20),.G_20_20(G_20),.P_21_21(P_21),.G_21_21(G_21),.P_22_22(P_22),.G_22_22(G_22),.P_23_23(P_23),.G_23_23(G_23),.P_24_24(P_24),.G_24_24(G_24),.P_25_25(P_25),.G_25_25(G_25),.P_26_26(P_26),.G_26_26(G_26),.P_27_27(P_27),.G_27_27(G_27),.P_28_28(P_28),.G_28_28(G_28),.P_29_29(P_29),.G_29_29(G_29),.P_30_30(P_30),.G_30_30(G_30),.P_31_31(P_31),.G_31_31(G_31),.P_32_32(P_32),.G_32_32(G_32),._P_0_0(P_0_0),._G_0_0(G_0_0),.P_1_0(P_1_0),.G_1_0(G_1_0),.P_2_0(P_2_0),.G_2_0(G_2_0),.P_3_0(P_3_0),.G_3_0(G_3_0),.P_4_0(P_4_0),.G_4_0(G_4_0),.P_5_0(P_5_0),.G_5_0(G_5_0),.P_6_0(P_6_0),.G_6_0(G_6_0),.P_7_0(P_7_0),.G_7_0(G_7_0),.P_8_0(P_8_0),.G_8_0(G_8_0),.P_9_0(P_9_0),.G_9_0(G_9_0),.P_10_0(P_10_0),.G_10_0(G_10_0),.P_11_0(P_11_0),.G_11_0(G_11_0),.P_12_0(P_12_0),.G_12_0(G_12_0),.P_13_0(P_13_0),.G_13_0(G_13_0),.P_14_0(P_14_0),.G_14_0(G_14_0),.P_15_0(P_15_0),.G_15_0(G_15_0),.P_16_0(P_16_0),.G_16_0(G_16_0),.P_17_0(P_17_0),.G_17_0(G_17_0),.P_18_0(P_18_0),.G_18_0(G_18_0),.P_19_0(P_19_0),.G_19_0(G_19_0),.P_20_0(P_20_0),.G_20_0(G_20_0),.P_21_0(P_21_0),.G_21_0(G_21_0),.P_22_0(P_22_0),.G_22_0(G_22_0),.P_23_0(P_23_0),.G_23_0(G_23_0),.P_24_0(P_24_0),.G_24_0(G_24_0),.P_25_0(P_25_0),.G_25_0(G_25_0),.P_26_0(P_26_0),.G_26_0(G_26_0),.P_27_0(P_27_0),.G_27_0(G_27_0),.P_28_0(P_28_0),.G_28_0(G_28_0),.P_29_0(P_29_0),.G_29_0(G_29_0),.P_30_0(P_30_0),.G_30_0(G_30_0),.P_31_0(P_31_0),.G_31_0(G_31_0),.P_32_0(P_32_0),.G_32_0(G_32_0));
SumLogic _SumLogic(.P_0(P_0),.G_0_0(G_0_0),.P_1(P_1),.G_1_0(G_1_0),.P_2(P_2),.G_2_0(G_2_0),.P_3(P_3),.G_3_0(G_3_0),.P_4(P_4),.G_4_0(G_4_0),.P_5(P_5),.G_5_0(G_5_0),.P_6(P_6),.G_6_0(G_6_0),.P_7(P_7),.G_7_0(G_7_0),.P_8(P_8),.G_8_0(G_8_0),.P_9(P_9),.G_9_0(G_9_0),.P_10(P_10),.G_10_0(G_10_0),.P_11(P_11),.G_11_0(G_11_0),.P_12(P_12),.G_12_0(G_12_0),.P_13(P_13),.G_13_0(G_13_0),.P_14(P_14),.G_14_0(G_14_0),.P_15(P_15),.G_15_0(G_15_0),.P_16(P_16),.G_16_0(G_16_0),.P_17(P_17),.G_17_0(G_17_0),.P_18(P_18),.G_18_0(G_18_0),.P_19(P_19),.G_19_0(G_19_0),.P_20(P_20),.G_20_0(G_20_0),.P_21(P_21),.G_21_0(G_21_0),.P_22(P_22),.G_22_0(G_22_0),.P_23(P_23),.G_23_0(G_23_0),.P_24(P_24),.G_24_0(G_24_0),.P_25(P_25),.G_25_0(G_25_0),.P_26(P_26),.G_26_0(G_26_0),.P_27(P_27),.G_27_0(G_27_0),.P_28(P_28),.G_28_0(G_28_0),.P_29(P_29),.G_29_0(G_29_0),.P_30(P_30),.G_30_0(G_30_0),.P_31(P_31),.G_31_0(G_31_0),.P_32(P_32),.G_32_0(G_32_0),.S_1(S_1),.S_2(S_2),.S_3(S_3),.S_4(S_4),.S_5(S_5),.S_6(S_6),.S_7(S_7),.S_8(S_8),.S_9(S_9),.S_10(S_10),.S_11(S_11),.S_12(S_12),.S_13(S_13),.S_14(S_14),.S_15(S_15),.S_16(S_16),.S_17(S_17),.S_18(S_18),.S_19(S_19),.S_20(S_20),.S_21(S_21),.S_22(S_22),.S_23(S_23),.S_24(S_24),.S_25(S_25),.S_26(S_26),.S_27(S_27),.S_28(S_28),.S_29(S_29),.S_30(S_30),.S_31(S_31),.S_32(S_32),.C_out(C_out));
endmodule
