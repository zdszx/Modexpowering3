module GroupPGLogic ( P_0_0,G_0_0,P_1_1,G_1_1,P_2_2,G_2_2,P_3_3,G_3_3,P_4_4,G_4_4,P_5_5,G_5_5,P_6_6,G_6_6,P_7_7,G_7_7,P_8_8,G_8_8,_P_0_0,_G_0_0,P_1_0,G_1_0,P_2_0,G_2_0,P_3_0,G_3_0,P_4_0,G_4_0,P_5_0,G_5_0,P_6_0,G_6_0,P_7_0,G_7_0,P_8_0,G_8_0 );
input P_0_0;
input G_0_0;
input P_1_1;
input G_1_1;
input P_2_2;
input G_2_2;
input P_3_3;
input G_3_3;
input P_4_4;
input G_4_4;
input P_5_5;
input G_5_5;
input P_6_6;
input G_6_6;
input P_7_7;
input G_7_7;
input P_8_8;
input G_8_8;
output _P_0_0;
output _G_0_0;
output P_1_0;
output G_1_0;
output P_2_0;
output G_2_0;
output P_3_0;
output G_3_0;
output P_4_0;
output G_4_0;
output P_5_0;
output G_5_0;
output P_6_0;
output G_6_0;
output P_7_0;
output G_7_0;
output P_8_0;
output G_8_0;
wire G_3_2;
wire P_3_2;
wire G_5_4;
wire P_5_4;
wire G_7_6;
wire P_7_6;
wire G_7_4;
wire P_7_4;
GrayBlock gray_block_1_0(.G_i_k(G_1_1),.P_i_k(P_1_1),.G_km1_j(G_0_0),.G_i_j(G_1_0));
BlackBlock black_block_3_2(.G_i_k(G_3_3),.P_i_k(P_3_3),.G_km1_j(G_2_2),.P_km1_j(P_2_2),.G_i_j(G_3_2),.P_i_j(P_3_2));
BlackBlock black_block_5_4(.G_i_k(G_5_5),.P_i_k(P_5_5),.G_km1_j(G_4_4),.P_km1_j(P_4_4),.G_i_j(G_5_4),.P_i_j(P_5_4));
BlackBlock black_block_7_6(.G_i_k(G_7_7),.P_i_k(P_7_7),.G_km1_j(G_6_6),.P_km1_j(P_6_6),.G_i_j(G_7_6),.P_i_j(P_7_6));
GrayBlock gray_block_3_0(.G_i_k(G_3_2),.P_i_k(P_3_2),.G_km1_j(G_1_0),.G_i_j(G_3_0));
BlackBlock black_block_7_4(.G_i_k(G_7_6),.P_i_k(P_7_6),.G_km1_j(G_5_4),.P_km1_j(P_5_4),.G_i_j(G_7_4),.P_i_j(P_7_4));
GrayBlock gray_block_7_0(.G_i_k(G_7_4),.P_i_k(P_7_4),.G_km1_j(G_3_0),.G_i_j(G_7_0));
GrayBlock gray_block_5_3(.G_i_k(G_5_4),.P_i_k(P_5_4),.G_km1_j(G_3_0),.G_i_j(G_5_0));
GrayBlock gray_block_2_1(.G_i_k(G_2_2),.P_i_k(P_2_2),.G_km1_j(G_1_0),.G_i_j(G_2_0));
GrayBlock gray_block_4_3(.G_i_k(G_4_4),.P_i_k(P_4_4),.G_km1_j(G_3_0),.G_i_j(G_4_0));
GrayBlock gray_block_6_5(.G_i_k(G_6_6),.P_i_k(P_6_6),.G_km1_j(G_5_0),.G_i_j(G_6_0));
GrayBlock gray_block_8_7(.G_i_k(G_8_8),.P_i_k(P_8_8),.G_km1_j(G_7_0),.G_i_j(G_8_0));
assign _P_0_0 = P_0_0 ;
assign _G_0_0 = G_0_0 ;
endmodule
