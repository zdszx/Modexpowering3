module test();
	reg[64:0] s_golden;
	reg[64:1] a,b;
	reg c_in;
	wire[64:1] s;

	BrentKungAdder adder(
							.A_1(a[1]), .B_1(b[1]),
							.A_2(a[2]), .B_2(b[2]),
							.A_3(a[3]), .B_3(b[3]),
							.A_4(a[4]), .B_4(b[4]),
							.A_5(a[5]), .B_5(b[5]),
							.A_6(a[6]), .B_6(b[6]),
							.A_7(a[7]), .B_7(b[7]),
							.A_8(a[8]), .B_8(b[8]),
							.A_9(a[9]), .B_9(b[9]),
							.A_10(a[10]), .B_10(b[10]),
							.A_11(a[11]), .B_11(b[11]),
							.A_12(a[12]), .B_12(b[12]),
							.A_13(a[13]), .B_13(b[13]),
							.A_14(a[14]), .B_14(b[14]),
							.A_15(a[15]), .B_15(b[15]),
							.A_16(a[16]), .B_16(b[16]),
							.A_17(a[17]), .B_17(b[17]),
							.A_18(a[18]), .B_18(b[18]),
							.A_19(a[19]), .B_19(b[19]),
							.A_20(a[20]), .B_20(b[20]),
							.A_21(a[21]), .B_21(b[21]),
							.A_22(a[22]), .B_22(b[22]),
							.A_23(a[23]), .B_23(b[23]),
							.A_24(a[24]), .B_24(b[24]),
							.A_25(a[25]), .B_25(b[25]),
							.A_26(a[26]), .B_26(b[26]),
							.A_27(a[27]), .B_27(b[27]),
							.A_28(a[28]), .B_28(b[28]),
							.A_29(a[29]), .B_29(b[29]),
							.A_30(a[30]), .B_30(b[30]),
							.A_31(a[31]), .B_31(b[31]),
							.A_32(a[32]), .B_32(b[32]),
							.A_33(a[33]), .B_33(b[33]),
							.A_34(a[34]), .B_34(b[34]),
							.A_35(a[35]), .B_35(b[35]),
							.A_36(a[36]), .B_36(b[36]),
							.A_37(a[37]), .B_37(b[37]),
							.A_38(a[38]), .B_38(b[38]),
							.A_39(a[39]), .B_39(b[39]),
							.A_40(a[40]), .B_40(b[40]),
							.A_41(a[41]), .B_41(b[41]),
							.A_42(a[42]), .B_42(b[42]),
							.A_43(a[43]), .B_43(b[43]),
							.A_44(a[44]), .B_44(b[44]),
							.A_45(a[45]), .B_45(b[45]),
							.A_46(a[46]), .B_46(b[46]),
							.A_47(a[47]), .B_47(b[47]),
							.A_48(a[48]), .B_48(b[48]),
							.A_49(a[49]), .B_49(b[49]),
							.A_50(a[50]), .B_50(b[50]),
							.A_51(a[51]), .B_51(b[51]),
							.A_52(a[52]), .B_52(b[52]),
							.A_53(a[53]), .B_53(b[53]),
							.A_54(a[54]), .B_54(b[54]),
							.A_55(a[55]), .B_55(b[55]),
							.A_56(a[56]), .B_56(b[56]),
							.A_57(a[57]), .B_57(b[57]),
							.A_58(a[58]), .B_58(b[58]),
							.A_59(a[59]), .B_59(b[59]),
							.A_60(a[60]), .B_60(b[60]),
							.A_61(a[61]), .B_61(b[61]),
							.A_62(a[62]), .B_62(b[62]),
							.A_63(a[63]), .B_63(b[63]),
							.A_64(a[64]), .B_64(b[64]),
							.C_0(c_in),
							.S_1(s[1]), .S_2(s[2]), 
							.S_3(s[3]), .S_4(s[4]), 
							.S_5(s[5]), .S_6(s[6]), 
							.S_7(s[7]), .S_8(s[8]), 
							.S_9(s[9]), .S_10(s[10]), 
							.S_11(s[11]), .S_12(s[12]), 
							.S_13(s[13]), .S_14(s[14]), 
							.S_15(s[15]), .S_16(s[16]), 
							.S_17(s[17]), .S_18(s[18]), 
							.S_19(s[19]), .S_20(s[20]), 
							.S_21(s[21]), .S_22(s[22]), 
							.S_23(s[23]), .S_24(s[24]), 
							.S_25(s[25]), .S_26(s[26]), 
							.S_27(s[27]), .S_28(s[28]), 
							.S_29(s[29]), .S_30(s[30]), 
							.S_31(s[31]), .S_32(s[32]), 
							.S_33(s[33]), .S_34(s[34]), 
							.S_35(s[35]), .S_36(s[36]), 
							.S_37(s[37]), .S_38(s[38]), 
							.S_39(s[39]), .S_40(s[40]), 
							.S_41(s[41]), .S_42(s[42]), 
							.S_43(s[43]), .S_44(s[44]), 
							.S_45(s[45]), .S_46(s[46]), 
							.S_47(s[47]), .S_48(s[48]), 
							.S_49(s[49]), .S_50(s[50]), 
							.S_51(s[51]), .S_52(s[52]), 
							.S_53(s[53]), .S_54(s[54]), 
							.S_55(s[55]), .S_56(s[56]), 
							.S_57(s[57]), .S_58(s[58]), 
							.S_59(s[59]), .S_60(s[60]), 
							.S_61(s[61]), .S_62(s[62]), 
							.S_63(s[63]), .S_64(s[64]), 
							.C_out(c_out));
	always @(a,b,c_in) begin
		s_golden = a + b + c_in;
	end

	initial begin
		c_in = 1'b0;
		a = 64'b00110011_00110011_00110011_00110011_00110011_00110011_00110011_00110011;
		b = 64'b00110011_00110011_00110011_00110011_00110011_00110011_00110011_00110001;
		#100
		$display("================================================================================================================");
		$display("In_1 = %d, In_2 = %d, c_in = %b, c_out = %b, My_Result = %d, Golden_Result = %d",a, b, c_in, c_out, s, s_golden);
		#100;
		c_in = 1'b0;
		a = 64'b10110011_00110011_00110011_00110011_00110011_00110011_00110011_00110101;
		b = 64'b10110011_00110011_00110011_00110011_00110011_00110011_00110011_00111100;
		#100
		$display("================================================================================================================");
		$display("In_1 = %d, In_2 = %d, c_in = %b, c_out = %b, My_Result = %d, Golden_Result = %d",a, b, c_in, c_out, s, s_golden);
		$display("================================================================================================================");
		#100;
	end
endmodule