module BitwisePGLogic ( A_1,B_1,A_2,B_2,A_3,B_3,A_4,B_4,A_5,B_5,A_6,B_6,A_7,B_7,A_8,B_8,A_9,B_9,A_10,B_10,A_11,B_11,A_12,B_12,A_13,B_13,A_14,B_14,A_15,B_15,A_16,B_16,A_17,B_17,A_18,B_18,A_19,B_19,A_20,B_20,A_21,B_21,A_22,B_22,A_23,B_23,A_24,B_24,A_25,B_25,A_26,B_26,A_27,B_27,A_28,B_28,A_29,B_29,A_30,B_30,A_31,B_31,A_32,B_32,A_33,B_33,A_34,B_34,A_35,B_35,A_36,B_36,A_37,B_37,A_38,B_38,A_39,B_39,A_40,B_40,A_41,B_41,A_42,B_42,A_43,B_43,A_44,B_44,A_45,B_45,A_46,B_46,A_47,B_47,A_48,B_48,A_49,B_49,A_50,B_50,A_51,B_51,A_52,B_52,A_53,B_53,A_54,B_54,A_55,B_55,A_56,B_56,A_57,B_57,A_58,B_58,A_59,B_59,A_60,B_60,A_61,B_61,A_62,B_62,A_63,B_63,A_64,B_64,C_0,P_0,G_0,P_1,G_1,P_2,G_2,P_3,G_3,P_4,G_4,P_5,G_5,P_6,G_6,P_7,G_7,P_8,G_8,P_9,G_9,P_10,G_10,P_11,G_11,P_12,G_12,P_13,G_13,P_14,G_14,P_15,G_15,P_16,G_16,P_17,G_17,P_18,G_18,P_19,G_19,P_20,G_20,P_21,G_21,P_22,G_22,P_23,G_23,P_24,G_24,P_25,G_25,P_26,G_26,P_27,G_27,P_28,G_28,P_29,G_29,P_30,G_30,P_31,G_31,P_32,G_32,P_33,G_33,P_34,G_34,P_35,G_35,P_36,G_36,P_37,G_37,P_38,G_38,P_39,G_39,P_40,G_40,P_41,G_41,P_42,G_42,P_43,G_43,P_44,G_44,P_45,G_45,P_46,G_46,P_47,G_47,P_48,G_48,P_49,G_49,P_50,G_50,P_51,G_51,P_52,G_52,P_53,G_53,P_54,G_54,P_55,G_55,P_56,G_56,P_57,G_57,P_58,G_58,P_59,G_59,P_60,G_60,P_61,G_61,P_62,G_62,P_63,G_63,P_64,G_64 );
input A_1;
input B_1;
input A_2;
input B_2;
input A_3;
input B_3;
input A_4;
input B_4;
input A_5;
input B_5;
input A_6;
input B_6;
input A_7;
input B_7;
input A_8;
input B_8;
input A_9;
input B_9;
input A_10;
input B_10;
input A_11;
input B_11;
input A_12;
input B_12;
input A_13;
input B_13;
input A_14;
input B_14;
input A_15;
input B_15;
input A_16;
input B_16;
input A_17;
input B_17;
input A_18;
input B_18;
input A_19;
input B_19;
input A_20;
input B_20;
input A_21;
input B_21;
input A_22;
input B_22;
input A_23;
input B_23;
input A_24;
input B_24;
input A_25;
input B_25;
input A_26;
input B_26;
input A_27;
input B_27;
input A_28;
input B_28;
input A_29;
input B_29;
input A_30;
input B_30;
input A_31;
input B_31;
input A_32;
input B_32;
input A_33;
input B_33;
input A_34;
input B_34;
input A_35;
input B_35;
input A_36;
input B_36;
input A_37;
input B_37;
input A_38;
input B_38;
input A_39;
input B_39;
input A_40;
input B_40;
input A_41;
input B_41;
input A_42;
input B_42;
input A_43;
input B_43;
input A_44;
input B_44;
input A_45;
input B_45;
input A_46;
input B_46;
input A_47;
input B_47;
input A_48;
input B_48;
input A_49;
input B_49;
input A_50;
input B_50;
input A_51;
input B_51;
input A_52;
input B_52;
input A_53;
input B_53;
input A_54;
input B_54;
input A_55;
input B_55;
input A_56;
input B_56;
input A_57;
input B_57;
input A_58;
input B_58;
input A_59;
input B_59;
input A_60;
input B_60;
input A_61;
input B_61;
input A_62;
input B_62;
input A_63;
input B_63;
input A_64;
input B_64;
input C_0;
output P_0;
output G_0;
output P_1;
output G_1;
output P_2;
output G_2;
output P_3;
output G_3;
output P_4;
output G_4;
output P_5;
output G_5;
output P_6;
output G_6;
output P_7;
output G_7;
output P_8;
output G_8;
output P_9;
output G_9;
output P_10;
output G_10;
output P_11;
output G_11;
output P_12;
output G_12;
output P_13;
output G_13;
output P_14;
output G_14;
output P_15;
output G_15;
output P_16;
output G_16;
output P_17;
output G_17;
output P_18;
output G_18;
output P_19;
output G_19;
output P_20;
output G_20;
output P_21;
output G_21;
output P_22;
output G_22;
output P_23;
output G_23;
output P_24;
output G_24;
output P_25;
output G_25;
output P_26;
output G_26;
output P_27;
output G_27;
output P_28;
output G_28;
output P_29;
output G_29;
output P_30;
output G_30;
output P_31;
output G_31;
output P_32;
output G_32;
output P_33;
output G_33;
output P_34;
output G_34;
output P_35;
output G_35;
output P_36;
output G_36;
output P_37;
output G_37;
output P_38;
output G_38;
output P_39;
output G_39;
output P_40;
output G_40;
output P_41;
output G_41;
output P_42;
output G_42;
output P_43;
output G_43;
output P_44;
output G_44;
output P_45;
output G_45;
output P_46;
output G_46;
output P_47;
output G_47;
output P_48;
output G_48;
output P_49;
output G_49;
output P_50;
output G_50;
output P_51;
output G_51;
output P_52;
output G_52;
output P_53;
output G_53;
output P_54;
output G_54;
output P_55;
output G_55;
output P_56;
output G_56;
output P_57;
output G_57;
output P_58;
output G_58;
output P_59;
output G_59;
output P_60;
output G_60;
output P_61;
output G_61;
output P_62;
output G_62;
output P_63;
output G_63;
output P_64;
output G_64;
// Bit 0
assign P_0 = 0 ;
assign G_0 = C_0 ;
// Bit 1
PG PG_Bit_1(.A_i(A_1),.B_i(B_1),.P_i(P_1),.G_i(G_1));
// Bit 2
PG PG_Bit_2(.A_i(A_2),.B_i(B_2),.P_i(P_2),.G_i(G_2));
// Bit 3
PG PG_Bit_3(.A_i(A_3),.B_i(B_3),.P_i(P_3),.G_i(G_3));
// Bit 4
PG PG_Bit_4(.A_i(A_4),.B_i(B_4),.P_i(P_4),.G_i(G_4));
// Bit 5
PG PG_Bit_5(.A_i(A_5),.B_i(B_5),.P_i(P_5),.G_i(G_5));
// Bit 6
PG PG_Bit_6(.A_i(A_6),.B_i(B_6),.P_i(P_6),.G_i(G_6));
// Bit 7
PG PG_Bit_7(.A_i(A_7),.B_i(B_7),.P_i(P_7),.G_i(G_7));
// Bit 8
PG PG_Bit_8(.A_i(A_8),.B_i(B_8),.P_i(P_8),.G_i(G_8));
// Bit 9
PG PG_Bit_9(.A_i(A_9),.B_i(B_9),.P_i(P_9),.G_i(G_9));
// Bit 10
PG PG_Bit_10(.A_i(A_10),.B_i(B_10),.P_i(P_10),.G_i(G_10));
// Bit 11
PG PG_Bit_11(.A_i(A_11),.B_i(B_11),.P_i(P_11),.G_i(G_11));
// Bit 12
PG PG_Bit_12(.A_i(A_12),.B_i(B_12),.P_i(P_12),.G_i(G_12));
// Bit 13
PG PG_Bit_13(.A_i(A_13),.B_i(B_13),.P_i(P_13),.G_i(G_13));
// Bit 14
PG PG_Bit_14(.A_i(A_14),.B_i(B_14),.P_i(P_14),.G_i(G_14));
// Bit 15
PG PG_Bit_15(.A_i(A_15),.B_i(B_15),.P_i(P_15),.G_i(G_15));
// Bit 16
PG PG_Bit_16(.A_i(A_16),.B_i(B_16),.P_i(P_16),.G_i(G_16));
// Bit 17
PG PG_Bit_17(.A_i(A_17),.B_i(B_17),.P_i(P_17),.G_i(G_17));
// Bit 18
PG PG_Bit_18(.A_i(A_18),.B_i(B_18),.P_i(P_18),.G_i(G_18));
// Bit 19
PG PG_Bit_19(.A_i(A_19),.B_i(B_19),.P_i(P_19),.G_i(G_19));
// Bit 20
PG PG_Bit_20(.A_i(A_20),.B_i(B_20),.P_i(P_20),.G_i(G_20));
// Bit 21
PG PG_Bit_21(.A_i(A_21),.B_i(B_21),.P_i(P_21),.G_i(G_21));
// Bit 22
PG PG_Bit_22(.A_i(A_22),.B_i(B_22),.P_i(P_22),.G_i(G_22));
// Bit 23
PG PG_Bit_23(.A_i(A_23),.B_i(B_23),.P_i(P_23),.G_i(G_23));
// Bit 24
PG PG_Bit_24(.A_i(A_24),.B_i(B_24),.P_i(P_24),.G_i(G_24));
// Bit 25
PG PG_Bit_25(.A_i(A_25),.B_i(B_25),.P_i(P_25),.G_i(G_25));
// Bit 26
PG PG_Bit_26(.A_i(A_26),.B_i(B_26),.P_i(P_26),.G_i(G_26));
// Bit 27
PG PG_Bit_27(.A_i(A_27),.B_i(B_27),.P_i(P_27),.G_i(G_27));
// Bit 28
PG PG_Bit_28(.A_i(A_28),.B_i(B_28),.P_i(P_28),.G_i(G_28));
// Bit 29
PG PG_Bit_29(.A_i(A_29),.B_i(B_29),.P_i(P_29),.G_i(G_29));
// Bit 30
PG PG_Bit_30(.A_i(A_30),.B_i(B_30),.P_i(P_30),.G_i(G_30));
// Bit 31
PG PG_Bit_31(.A_i(A_31),.B_i(B_31),.P_i(P_31),.G_i(G_31));
// Bit 32
PG PG_Bit_32(.A_i(A_32),.B_i(B_32),.P_i(P_32),.G_i(G_32));
// Bit 33
PG PG_Bit_33(.A_i(A_33),.B_i(B_33),.P_i(P_33),.G_i(G_33));
// Bit 34
PG PG_Bit_34(.A_i(A_34),.B_i(B_34),.P_i(P_34),.G_i(G_34));
// Bit 35
PG PG_Bit_35(.A_i(A_35),.B_i(B_35),.P_i(P_35),.G_i(G_35));
// Bit 36
PG PG_Bit_36(.A_i(A_36),.B_i(B_36),.P_i(P_36),.G_i(G_36));
// Bit 37
PG PG_Bit_37(.A_i(A_37),.B_i(B_37),.P_i(P_37),.G_i(G_37));
// Bit 38
PG PG_Bit_38(.A_i(A_38),.B_i(B_38),.P_i(P_38),.G_i(G_38));
// Bit 39
PG PG_Bit_39(.A_i(A_39),.B_i(B_39),.P_i(P_39),.G_i(G_39));
// Bit 40
PG PG_Bit_40(.A_i(A_40),.B_i(B_40),.P_i(P_40),.G_i(G_40));
// Bit 41
PG PG_Bit_41(.A_i(A_41),.B_i(B_41),.P_i(P_41),.G_i(G_41));
// Bit 42
PG PG_Bit_42(.A_i(A_42),.B_i(B_42),.P_i(P_42),.G_i(G_42));
// Bit 43
PG PG_Bit_43(.A_i(A_43),.B_i(B_43),.P_i(P_43),.G_i(G_43));
// Bit 44
PG PG_Bit_44(.A_i(A_44),.B_i(B_44),.P_i(P_44),.G_i(G_44));
// Bit 45
PG PG_Bit_45(.A_i(A_45),.B_i(B_45),.P_i(P_45),.G_i(G_45));
// Bit 46
PG PG_Bit_46(.A_i(A_46),.B_i(B_46),.P_i(P_46),.G_i(G_46));
// Bit 47
PG PG_Bit_47(.A_i(A_47),.B_i(B_47),.P_i(P_47),.G_i(G_47));
// Bit 48
PG PG_Bit_48(.A_i(A_48),.B_i(B_48),.P_i(P_48),.G_i(G_48));
// Bit 49
PG PG_Bit_49(.A_i(A_49),.B_i(B_49),.P_i(P_49),.G_i(G_49));
// Bit 50
PG PG_Bit_50(.A_i(A_50),.B_i(B_50),.P_i(P_50),.G_i(G_50));
// Bit 51
PG PG_Bit_51(.A_i(A_51),.B_i(B_51),.P_i(P_51),.G_i(G_51));
// Bit 52
PG PG_Bit_52(.A_i(A_52),.B_i(B_52),.P_i(P_52),.G_i(G_52));
// Bit 53
PG PG_Bit_53(.A_i(A_53),.B_i(B_53),.P_i(P_53),.G_i(G_53));
// Bit 54
PG PG_Bit_54(.A_i(A_54),.B_i(B_54),.P_i(P_54),.G_i(G_54));
// Bit 55
PG PG_Bit_55(.A_i(A_55),.B_i(B_55),.P_i(P_55),.G_i(G_55));
// Bit 56
PG PG_Bit_56(.A_i(A_56),.B_i(B_56),.P_i(P_56),.G_i(G_56));
// Bit 57
PG PG_Bit_57(.A_i(A_57),.B_i(B_57),.P_i(P_57),.G_i(G_57));
// Bit 58
PG PG_Bit_58(.A_i(A_58),.B_i(B_58),.P_i(P_58),.G_i(G_58));
// Bit 59
PG PG_Bit_59(.A_i(A_59),.B_i(B_59),.P_i(P_59),.G_i(G_59));
// Bit 60
PG PG_Bit_60(.A_i(A_60),.B_i(B_60),.P_i(P_60),.G_i(G_60));
// Bit 61
PG PG_Bit_61(.A_i(A_61),.B_i(B_61),.P_i(P_61),.G_i(G_61));
// Bit 62
PG PG_Bit_62(.A_i(A_62),.B_i(B_62),.P_i(P_62),.G_i(G_62));
// Bit 63
PG PG_Bit_63(.A_i(A_63),.B_i(B_63),.P_i(P_63),.G_i(G_63));
// Bit 64
PG PG_Bit_64(.A_i(A_64),.B_i(B_64),.P_i(P_64),.G_i(G_64));
endmodule
