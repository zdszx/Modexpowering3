module BrentKungAdder ( A_1,B_1,A_2,B_2,A_3,B_3,A_4,B_4,C_0,S_1,S_2,S_3,S_4,C_out );
input A_1;
input B_1;
input A_2;
input B_2;
input A_3;
input B_3;
input A_4;
input B_4;
input C_0;
output S_1;
output S_2;
output S_3;
output S_4;
output C_out;
wire P_0;
wire G_0;
wire P_1;
wire G_1;
wire P_2;
wire G_2;
wire P_3;
wire G_3;
wire P_4;
wire G_4;
wire P_0_0;
wire G_0_0;
wire P_1_0;
wire G_1_0;
wire P_2_0;
wire G_2_0;
wire P_3_0;
wire G_3_0;
wire P_4_0;
wire G_4_0;
BitwisePGLogic _BitwisePGLogic(.C_0(C_0),.A_1(A_1),.B_1(B_1),.A_2(A_2),.B_2(B_2),.A_3(A_3),.B_3(B_3),.A_4(A_4),.B_4(B_4),.P_0(P_0),.G_0(G_0),.P_1(P_1),.G_1(G_1),.P_2(P_2),.G_2(G_2),.P_3(P_3),.G_3(G_3),.P_4(P_4),.G_4(G_4));
GroupPGLogic _GroupPGLogic(.P_0_0(P_0),.G_0_0(G_0),.P_1_1(P_1),.G_1_1(G_1),.P_2_2(P_2),.G_2_2(G_2),.P_3_3(P_3),.G_3_3(G_3),.P_4_4(P_4),.G_4_4(G_4),._P_0_0(P_0_0),._G_0_0(G_0_0),.P_1_0(P_1_0),.G_1_0(G_1_0),.P_2_0(P_2_0),.G_2_0(G_2_0),.P_3_0(P_3_0),.G_3_0(G_3_0),.P_4_0(P_4_0),.G_4_0(G_4_0));
SumLogic _SumLogic(.P_0(P_0),.G_0_0(G_0_0),.P_1(P_1),.G_1_0(G_1_0),.P_2(P_2),.G_2_0(G_2_0),.P_3(P_3),.G_3_0(G_3_0),.P_4(P_4),.G_4_0(G_4_0),.S_1(S_1),.S_2(S_2),.S_3(S_3),.S_4(S_4),.C_out(C_out));
endmodule
