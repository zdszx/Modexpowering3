module test();
	reg[32:0] s_golden;
	reg[32:1] a,b;
	reg c_in;
	wire[32:1] s;

	BrentKungAdder adder(
							.A_1(a[1]), .B_1(b[1]),
							.A_2(a[2]), .B_2(b[2]),
							.A_3(a[3]), .B_3(b[3]),
							.A_4(a[4]), .B_4(b[4]),
							.A_5(a[5]), .B_5(b[5]),
							.A_6(a[6]), .B_6(b[6]),
							.A_7(a[7]), .B_7(b[7]),
							.A_8(a[8]), .B_8(b[8]),
							.A_9(a[9]), .B_9(b[9]),
							.A_10(a[10]), .B_10(b[10]),
							.A_11(a[11]), .B_11(b[11]),
							.A_12(a[12]), .B_12(b[12]),
							.A_13(a[13]), .B_13(b[13]),
							.A_14(a[14]), .B_14(b[14]),
							.A_15(a[15]), .B_15(b[15]),
							.A_16(a[16]), .B_16(b[16]),
							.A_17(a[17]), .B_17(b[17]),
							.A_18(a[18]), .B_18(b[18]),
							.A_19(a[19]), .B_19(b[19]),
							.A_20(a[20]), .B_20(b[20]),
							.A_21(a[21]), .B_21(b[21]),
							.A_22(a[22]), .B_22(b[22]),
							.A_23(a[23]), .B_23(b[23]),
							.A_24(a[24]), .B_24(b[24]),
							.A_25(a[25]), .B_25(b[25]),
							.A_26(a[26]), .B_26(b[26]),
							.A_27(a[27]), .B_27(b[27]),
							.A_28(a[28]), .B_28(b[28]),
							.A_29(a[29]), .B_29(b[29]),
							.A_30(a[30]), .B_30(b[30]),
							.A_31(a[31]), .B_31(b[31]),
							.A_32(a[32]), .B_32(b[32]),
							.C_0(c_in),
							.S_1(s[1]), .S_2(s[2]), 
							.S_3(s[3]), .S_4(s[4]), 
							.S_5(s[5]), .S_6(s[6]), 
							.S_7(s[7]), .S_8(s[8]), 
							.S_9(s[9]), .S_10(s[10]), 
							.S_11(s[11]), .S_12(s[12]), 
							.S_13(s[13]), .S_14(s[14]), 
							.S_15(s[15]), .S_16(s[16]), 
							.S_17(s[17]), .S_18(s[18]), 
							.S_19(s[19]), .S_20(s[20]), 
							.S_21(s[21]), .S_22(s[22]), 
							.S_23(s[23]), .S_24(s[24]), 
							.S_25(s[25]), .S_26(s[26]), 
							.S_27(s[27]), .S_28(s[28]), 
							.S_29(s[29]), .S_30(s[30]), 
							.S_31(s[31]), .S_32(s[32]), 
							.C_out(c_out));
	always @(a,b,c_in) begin
		s_golden = a + b + c_in;
	end

	initial begin
		c_in = 1'b0;
		a = 32'b1000_1000_1011_0011_1000_1000_1011_0011;
		b = 32'b1000_1000_1011_0001_1000_1000_1011_0001;
		#100
		$display("================================================================================================================");
		$display("In_1 = %d, In_2 = %d, c_in = %b, c_out = %b, My_Result = %d, Golden_Result = %d",a, b, c_in, c_out, s, s_golden);
		#100;
		c_in = 1'b0;
		a = 32'b10000101;
		b = 32'b10001100;
		#100
		$display("================================================================================================================");
		$display("In_1 = %d, In_2 = %d, c_in = %b, c_out = %b, My_Result = %d, Golden_Result = %d",a, b, c_in, c_out, s, s_golden);
		$display("================================================================================================================");
		#100;
	end
endmodule